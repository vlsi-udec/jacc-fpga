`timescale 1ns / 1ps

module mmh3_f64 (
	input logic [0:0] clk,
	output logic [63:0] hash,
	input logic [61:0] in_data,
	input logic [0:0] in_valid,
	output logic [0:0] out_valid
);

logic [63:0] k[7:0];
logic [63:0] tmp[2:0];
logic [31:0] k1_m[9:0];
logic [32:0] k1_t0[5:0];
logic [33:0] k1_t1[3:0];
logic [63:0] k1_t2[1:0];
logic [63:0] k1_b[3:0];
logic [31:0] k4_m[9:0];
logic [32:0] k4_t0[5:0];
logic [33:0] k4_t1[3:0];
logic [63:0] k4_t2[1:0];
logic [63:0] k4_b[3:0];
logic [17:0] in_valid_r = 18'd0;

always_ff @(posedge clk) begin
	k[0] <= in_data >> 6'd33;
	tmp[0] <= in_data;
	k[1] <= tmp[0] ^ k[0];
	k1_b[0] <= k[1];
	k1_b[1] <= k[1];
	k1_b[2] <= k[1];
	k1_b[3] <= k[1];
	k1_m[0] <= k1_b[0][15:0] * 16'd36045;
	k1_m[1] <= k1_b[0][31:16] * 16'd36045;
	k1_m[2] <= k1_b[0][47:32] * 16'd36045;
	k1_m[3] <= k1_b[0][63:48] * 16'd36045;
	k1_m[4] <= k1_b[1][15:0] * 16'd60757;
	k1_m[5] <= k1_b[1][31:16] * 16'd60757;
	k1_m[6] <= k1_b[1][47:32] * 16'd60757;
	k1_m[7] <= k1_b[2][15:0] * 16'd45015;
	k1_m[8] <= k1_b[2][31:16] * 16'd45015;
	k1_m[9] <= k1_b[3][15:0] * 16'd65361;
	k1_t0[0] <= k1_m[0];
	k1_t0[1] <= k1_m[1] + k1_m[4];
	k1_t0[2] <= k1_m[2] + k1_m[5];
	k1_t0[3] <= k1_m[7];
	k1_t0[4] <= k1_m[3] + k1_m[6];
	k1_t0[5] <= k1_m[8] + k1_m[9];
	k1_t1[0] <= k1_t0[0];
	k1_t1[1] <= k1_t0[1];
	k1_t1[2] <= k1_t0[2] + k1_t0[3];
	k1_t1[3] <= k1_t0[4] + k1_t0[5];
	k1_t2[0] <= k1_t1[0] + (k1_t1[1] << 5'd16);
	k1_t2[1] <= k1_t1[2] + (k1_t1[3] << 5'd16);
	k[2] <= k1_t2[0] + (k1_t2[1] << 6'd32);
	k[3] <= k[2] >> 6'd33;
	tmp[1] <= k[2];
	k[4] <= tmp[1] ^ k[3];
	k4_b[0] <= k[4];
	k4_b[1] <= k[4];
	k4_b[2] <= k[4];
	k4_b[3] <= k[4];
	k4_m[0] <= k4_b[0][15:0] * 16'd60499;
	k4_m[1] <= k4_b[0][31:16] * 16'd60499;
	k4_m[2] <= k4_b[0][47:32] * 16'd60499;
	k4_m[3] <= k4_b[0][63:48] * 16'd60499;
	k4_m[4] <= k4_b[1][15:0] * 16'd6789;
	k4_m[5] <= k4_b[1][31:16] * 16'd6789;
	k4_m[6] <= k4_b[1][47:32] * 16'd6789;
	k4_m[7] <= k4_b[2][15:0] * 16'd47614;
	k4_m[8] <= k4_b[2][31:16] * 16'd47614;
	k4_m[9] <= k4_b[3][15:0] * 16'd50382;
	k4_t0[0] <= k4_m[0];
	k4_t0[1] <= k4_m[1] + k4_m[4];
	k4_t0[2] <= k4_m[2] + k4_m[5];
	k4_t0[3] <= k4_m[7];
	k4_t0[4] <= k4_m[3] + k4_m[6];
	k4_t0[5] <= k4_m[8] + k4_m[9];
	k4_t1[0] <= k4_t0[0];
	k4_t1[1] <= k4_t0[1];
	k4_t1[2] <= k4_t0[2] + k4_t0[3];
	k4_t1[3] <= k4_t0[4] + k4_t0[5];
	k4_t2[0] <= k4_t1[0] + (k4_t1[1] << 5'd16);
	k4_t2[1] <= k4_t1[2] + (k4_t1[3] << 5'd16);
	k[5] <= k4_t2[0] + (k4_t2[1] << 6'd32);
	k[6] <= k[5] >> 6'd33;
	tmp[2] <= k[5];
	k[7] <= tmp[2] ^ k[6];
	in_valid_r <= {in_valid_r[16:0], in_valid};
end

always_comb begin
	hash = k[7];
	out_valid = in_valid_r[17];
end

endmodule

