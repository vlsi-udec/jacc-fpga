`timescale 1ns / 1ps

module krnl_card_rtl (
	input wire [0:0] ap_clk,
	input wire [0:0] ap_clk_2,
	input wire [0:0] ap_rst_n,
	input wire [0:0] ap_rst_n_2,
	output wire [63:0] m_axi_gmem_ARADDR,
	output wire [1:0] m_axi_gmem_ARBURST,
	output wire [3:0] m_axi_gmem_ARCACHE,
	output wire [0:0] m_axi_gmem_ARID,
	output wire [7:0] m_axi_gmem_ARLEN,
	output wire [1:0] m_axi_gmem_ARLOCK,
	output wire [2:0] m_axi_gmem_ARPROT,
	output wire [3:0] m_axi_gmem_ARQOS,
	input wire [0:0] m_axi_gmem_ARREADY,
	output wire [3:0] m_axi_gmem_ARREGION,
	output wire [2:0] m_axi_gmem_ARSIZE,
	output wire [0:0] m_axi_gmem_ARVALID,
	output wire [63:0] m_axi_gmem_AWADDR,
	output wire [1:0] m_axi_gmem_AWBURST,
	output wire [3:0] m_axi_gmem_AWCACHE,
	output wire [0:0] m_axi_gmem_AWID,
	output wire [7:0] m_axi_gmem_AWLEN,
	output wire [1:0] m_axi_gmem_AWLOCK,
	output wire [2:0] m_axi_gmem_AWPROT,
	output wire [3:0] m_axi_gmem_AWQOS,
	input wire [0:0] m_axi_gmem_AWREADY,
	output wire [3:0] m_axi_gmem_AWREGION,
	output wire [2:0] m_axi_gmem_AWSIZE,
	output wire [0:0] m_axi_gmem_AWVALID,
	input wire [0:0] m_axi_gmem_BID,
	output wire [0:0] m_axi_gmem_BREADY,
	input wire [1:0] m_axi_gmem_BRESP,
	input wire [0:0] m_axi_gmem_BVALID,
	input wire [63:0] m_axi_gmem_RDATA,
	input wire [0:0] m_axi_gmem_RID,
	input wire [0:0] m_axi_gmem_RLAST,
	output wire [0:0] m_axi_gmem_RREADY,
	input wire [1:0] m_axi_gmem_RRESP,
	input wire [0:0] m_axi_gmem_RVALID,
	output wire [63:0] m_axi_gmem_WDATA,
	output wire [0:0] m_axi_gmem_WLAST,
	input wire [0:0] m_axi_gmem_WREADY,
	output wire [7:0] m_axi_gmem_WSTRB,
	output wire [0:0] m_axi_gmem_WVALID,
	input wire [63:0] p0_TDATA,
	output wire [0:0] p0_TREADY,
	input wire [0:0] p0_TVALID,
	input wire [63:0] p1_TDATA,
	output wire [0:0] p1_TREADY,
	input wire [0:0] p1_TVALID,
	input wire [63:0] p2_TDATA,
	output wire [0:0] p2_TREADY,
	input wire [0:0] p2_TVALID,
	input wire [63:0] p3_TDATA,
	output wire [0:0] p3_TREADY,
	input wire [0:0] p3_TVALID,
	input wire [63:0] p4_TDATA,
	output wire [0:0] p4_TREADY,
	input wire [0:0] p4_TVALID,
	input wire [63:0] p5_TDATA,
	output wire [0:0] p5_TREADY,
	input wire [0:0] p5_TVALID,
	input wire [63:0] p6_TDATA,
	output wire [0:0] p6_TREADY,
	input wire [0:0] p6_TVALID,
	input wire [63:0] p7_TDATA,
	output wire [0:0] p7_TREADY,
	input wire [0:0] p7_TVALID,
	input wire [31:0] s_axi_control_ARADDR,
	output wire [0:0] s_axi_control_ARREADY,
	input wire [0:0] s_axi_control_ARVALID,
	input wire [31:0] s_axi_control_AWADDR,
	output wire [0:0] s_axi_control_AWREADY,
	input wire [0:0] s_axi_control_AWVALID,
	input wire [0:0] s_axi_control_BREADY,
	output wire [1:0] s_axi_control_BRESP,
	output wire [0:0] s_axi_control_BVALID,
	output wire [31:0] s_axi_control_RDATA,
	input wire [0:0] s_axi_control_RREADY,
	output wire [1:0] s_axi_control_RRESP,
	output wire [0:0] s_axi_control_RVALID,
	input wire [31:0] s_axi_control_WDATA,
	output wire [0:0] s_axi_control_WREADY,
	input wire [3:0] s_axi_control_WSTRB,
	input wire [0:0] s_axi_control_WVALID
);


krnl_card_rtl_int krnl_card_rtl_int_inst0 (
	.ap_aclk (ap_clk),
	.ap_aclk_2 (ap_clk_2),
	.ap_rst_n (ap_rst_n),
	.ap_rst_n_2 (ap_rst_n_2),
	.m_axi_gmem_ARADDR (m_axi_gmem_ARADDR),
	.m_axi_gmem_ARBURST (m_axi_gmem_ARBURST),
	.m_axi_gmem_ARCACHE (m_axi_gmem_ARCACHE),
	.m_axi_gmem_ARID (m_axi_gmem_ARID),
	.m_axi_gmem_ARLEN (m_axi_gmem_ARLEN),
	.m_axi_gmem_ARLOCK (m_axi_gmem_ARLOCK),
	.m_axi_gmem_ARPROT (m_axi_gmem_ARPROT),
	.m_axi_gmem_ARQOS (m_axi_gmem_ARQOS),
	.m_axi_gmem_ARREADY (m_axi_gmem_ARREADY),
	.m_axi_gmem_ARREGION (m_axi_gmem_ARREGION),
	.m_axi_gmem_ARSIZE (m_axi_gmem_ARSIZE),
	.m_axi_gmem_ARVALID (m_axi_gmem_ARVALID),
	.m_axi_gmem_AWADDR (m_axi_gmem_AWADDR),
	.m_axi_gmem_AWBURST (m_axi_gmem_AWBURST),
	.m_axi_gmem_AWCACHE (m_axi_gmem_AWCACHE),
	.m_axi_gmem_AWID (m_axi_gmem_AWID),
	.m_axi_gmem_AWLEN (m_axi_gmem_AWLEN),
	.m_axi_gmem_AWLOCK (m_axi_gmem_AWLOCK),
	.m_axi_gmem_AWPROT (m_axi_gmem_AWPROT),
	.m_axi_gmem_AWQOS (m_axi_gmem_AWQOS),
	.m_axi_gmem_AWREADY (m_axi_gmem_AWREADY),
	.m_axi_gmem_AWREGION (m_axi_gmem_AWREGION),
	.m_axi_gmem_AWSIZE (m_axi_gmem_AWSIZE),
	.m_axi_gmem_AWVALID (m_axi_gmem_AWVALID),
	.m_axi_gmem_BID (m_axi_gmem_BID),
	.m_axi_gmem_BREADY (m_axi_gmem_BREADY),
	.m_axi_gmem_BRESP (m_axi_gmem_BRESP),
	.m_axi_gmem_BVALID (m_axi_gmem_BVALID),
	.m_axi_gmem_RDATA (m_axi_gmem_RDATA),
	.m_axi_gmem_RID (m_axi_gmem_RID),
	.m_axi_gmem_RLAST (m_axi_gmem_RLAST),
	.m_axi_gmem_RREADY (m_axi_gmem_RREADY),
	.m_axi_gmem_RRESP (m_axi_gmem_RRESP),
	.m_axi_gmem_RVALID (m_axi_gmem_RVALID),
	.m_axi_gmem_WDATA (m_axi_gmem_WDATA),
	.m_axi_gmem_WLAST (m_axi_gmem_WLAST),
	.m_axi_gmem_WREADY (m_axi_gmem_WREADY),
	.m_axi_gmem_WSTRB (m_axi_gmem_WSTRB),
	.m_axi_gmem_WVALID (m_axi_gmem_WVALID),
	.p0_TDATA (p0_TDATA),
	.p0_TREADY (p0_TREADY),
	.p0_TVALID (p0_TVALID),
	.p1_TDATA (p1_TDATA),
	.p1_TREADY (p1_TREADY),
	.p1_TVALID (p1_TVALID),
	.p2_TDATA (p2_TDATA),
	.p2_TREADY (p2_TREADY),
	.p2_TVALID (p2_TVALID),
	.p3_TDATA (p3_TDATA),
	.p3_TREADY (p3_TREADY),
	.p3_TVALID (p3_TVALID),
	.p4_TDATA (p4_TDATA),
	.p4_TREADY (p4_TREADY),
	.p4_TVALID (p4_TVALID),
	.p5_TDATA (p5_TDATA),
	.p5_TREADY (p5_TREADY),
	.p5_TVALID (p5_TVALID),
	.p6_TDATA (p6_TDATA),
	.p6_TREADY (p6_TREADY),
	.p6_TVALID (p6_TVALID),
	.p7_TDATA (p7_TDATA),
	.p7_TREADY (p7_TREADY),
	.p7_TVALID (p7_TVALID),
	.s_axi_control_ARADDR (s_axi_control_ARADDR),
	.s_axi_control_ARREADY (s_axi_control_ARREADY),
	.s_axi_control_ARVALID (s_axi_control_ARVALID),
	.s_axi_control_AWADDR (s_axi_control_AWADDR),
	.s_axi_control_AWREADY (s_axi_control_AWREADY),
	.s_axi_control_AWVALID (s_axi_control_AWVALID),
	.s_axi_control_BREADY (s_axi_control_BREADY),
	.s_axi_control_BRESP (s_axi_control_BRESP),
	.s_axi_control_BVALID (s_axi_control_BVALID),
	.s_axi_control_RDATA (s_axi_control_RDATA),
	.s_axi_control_RREADY (s_axi_control_RREADY),
	.s_axi_control_RRESP (s_axi_control_RRESP),
	.s_axi_control_RVALID (s_axi_control_RVALID),
	.s_axi_control_WDATA (s_axi_control_WDATA),
	.s_axi_control_WREADY (s_axi_control_WREADY),
	.s_axi_control_WSTRB (s_axi_control_WSTRB),
	.s_axi_control_WVALID (s_axi_control_WVALID)
);

endmodule

