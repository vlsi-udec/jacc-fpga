`timescale 1ns / 1ps

module krnl_hll_rtl (
	input wire [0:0] ap_clk,
	input wire [0:0] ap_clk_2,
	input wire [0:0] ap_rst_n,
	input wire [0:0] ap_rst_n_2,
	output wire [63:0] m_axi_gmem_0_ARADDR,
	output wire [1:0] m_axi_gmem_0_ARBURST,
	output wire [3:0] m_axi_gmem_0_ARCACHE,
	output wire [0:0] m_axi_gmem_0_ARID,
	output wire [7:0] m_axi_gmem_0_ARLEN,
	output wire [1:0] m_axi_gmem_0_ARLOCK,
	output wire [2:0] m_axi_gmem_0_ARPROT,
	output wire [3:0] m_axi_gmem_0_ARQOS,
	input wire [0:0] m_axi_gmem_0_ARREADY,
	output wire [3:0] m_axi_gmem_0_ARREGION,
	output wire [2:0] m_axi_gmem_0_ARSIZE,
	output wire [0:0] m_axi_gmem_0_ARVALID,
	output wire [63:0] m_axi_gmem_0_AWADDR,
	output wire [1:0] m_axi_gmem_0_AWBURST,
	output wire [3:0] m_axi_gmem_0_AWCACHE,
	output wire [0:0] m_axi_gmem_0_AWID,
	output wire [7:0] m_axi_gmem_0_AWLEN,
	output wire [1:0] m_axi_gmem_0_AWLOCK,
	output wire [2:0] m_axi_gmem_0_AWPROT,
	output wire [3:0] m_axi_gmem_0_AWQOS,
	input wire [0:0] m_axi_gmem_0_AWREADY,
	output wire [3:0] m_axi_gmem_0_AWREGION,
	output wire [2:0] m_axi_gmem_0_AWSIZE,
	output wire [0:0] m_axi_gmem_0_AWVALID,
	input wire [0:0] m_axi_gmem_0_BID,
	output wire [0:0] m_axi_gmem_0_BREADY,
	input wire [1:0] m_axi_gmem_0_BRESP,
	input wire [0:0] m_axi_gmem_0_BVALID,
	input wire [511:0] m_axi_gmem_0_RDATA,
	input wire [0:0] m_axi_gmem_0_RID,
	input wire [0:0] m_axi_gmem_0_RLAST,
	output wire [0:0] m_axi_gmem_0_RREADY,
	input wire [1:0] m_axi_gmem_0_RRESP,
	input wire [0:0] m_axi_gmem_0_RVALID,
	output wire [511:0] m_axi_gmem_0_WDATA,
	output wire [0:0] m_axi_gmem_0_WLAST,
	input wire [0:0] m_axi_gmem_0_WREADY,
	output wire [63:0] m_axi_gmem_0_WSTRB,
	output wire [0:0] m_axi_gmem_0_WVALID,
	output wire [63:0] m_axi_gmem_1_ARADDR,
	output wire [1:0] m_axi_gmem_1_ARBURST,
	output wire [3:0] m_axi_gmem_1_ARCACHE,
	output wire [0:0] m_axi_gmem_1_ARID,
	output wire [7:0] m_axi_gmem_1_ARLEN,
	output wire [1:0] m_axi_gmem_1_ARLOCK,
	output wire [2:0] m_axi_gmem_1_ARPROT,
	output wire [3:0] m_axi_gmem_1_ARQOS,
	input wire [0:0] m_axi_gmem_1_ARREADY,
	output wire [3:0] m_axi_gmem_1_ARREGION,
	output wire [2:0] m_axi_gmem_1_ARSIZE,
	output wire [0:0] m_axi_gmem_1_ARVALID,
	output wire [63:0] m_axi_gmem_1_AWADDR,
	output wire [1:0] m_axi_gmem_1_AWBURST,
	output wire [3:0] m_axi_gmem_1_AWCACHE,
	output wire [0:0] m_axi_gmem_1_AWID,
	output wire [7:0] m_axi_gmem_1_AWLEN,
	output wire [1:0] m_axi_gmem_1_AWLOCK,
	output wire [2:0] m_axi_gmem_1_AWPROT,
	output wire [3:0] m_axi_gmem_1_AWQOS,
	input wire [0:0] m_axi_gmem_1_AWREADY,
	output wire [3:0] m_axi_gmem_1_AWREGION,
	output wire [2:0] m_axi_gmem_1_AWSIZE,
	output wire [0:0] m_axi_gmem_1_AWVALID,
	input wire [0:0] m_axi_gmem_1_BID,
	output wire [0:0] m_axi_gmem_1_BREADY,
	input wire [1:0] m_axi_gmem_1_BRESP,
	input wire [0:0] m_axi_gmem_1_BVALID,
	input wire [511:0] m_axi_gmem_1_RDATA,
	input wire [0:0] m_axi_gmem_1_RID,
	input wire [0:0] m_axi_gmem_1_RLAST,
	output wire [0:0] m_axi_gmem_1_RREADY,
	input wire [1:0] m_axi_gmem_1_RRESP,
	input wire [0:0] m_axi_gmem_1_RVALID,
	output wire [511:0] m_axi_gmem_1_WDATA,
	output wire [0:0] m_axi_gmem_1_WLAST,
	input wire [0:0] m_axi_gmem_1_WREADY,
	output wire [63:0] m_axi_gmem_1_WSTRB,
	output wire [0:0] m_axi_gmem_1_WVALID,
	output wire [63:0] m_axi_gmem_2_ARADDR,
	output wire [1:0] m_axi_gmem_2_ARBURST,
	output wire [3:0] m_axi_gmem_2_ARCACHE,
	output wire [0:0] m_axi_gmem_2_ARID,
	output wire [7:0] m_axi_gmem_2_ARLEN,
	output wire [1:0] m_axi_gmem_2_ARLOCK,
	output wire [2:0] m_axi_gmem_2_ARPROT,
	output wire [3:0] m_axi_gmem_2_ARQOS,
	input wire [0:0] m_axi_gmem_2_ARREADY,
	output wire [3:0] m_axi_gmem_2_ARREGION,
	output wire [2:0] m_axi_gmem_2_ARSIZE,
	output wire [0:0] m_axi_gmem_2_ARVALID,
	output wire [63:0] m_axi_gmem_2_AWADDR,
	output wire [1:0] m_axi_gmem_2_AWBURST,
	output wire [3:0] m_axi_gmem_2_AWCACHE,
	output wire [0:0] m_axi_gmem_2_AWID,
	output wire [7:0] m_axi_gmem_2_AWLEN,
	output wire [1:0] m_axi_gmem_2_AWLOCK,
	output wire [2:0] m_axi_gmem_2_AWPROT,
	output wire [3:0] m_axi_gmem_2_AWQOS,
	input wire [0:0] m_axi_gmem_2_AWREADY,
	output wire [3:0] m_axi_gmem_2_AWREGION,
	output wire [2:0] m_axi_gmem_2_AWSIZE,
	output wire [0:0] m_axi_gmem_2_AWVALID,
	input wire [0:0] m_axi_gmem_2_BID,
	output wire [0:0] m_axi_gmem_2_BREADY,
	input wire [1:0] m_axi_gmem_2_BRESP,
	input wire [0:0] m_axi_gmem_2_BVALID,
	input wire [511:0] m_axi_gmem_2_RDATA,
	input wire [0:0] m_axi_gmem_2_RID,
	input wire [0:0] m_axi_gmem_2_RLAST,
	output wire [0:0] m_axi_gmem_2_RREADY,
	input wire [1:0] m_axi_gmem_2_RRESP,
	input wire [0:0] m_axi_gmem_2_RVALID,
	output wire [511:0] m_axi_gmem_2_WDATA,
	output wire [0:0] m_axi_gmem_2_WLAST,
	input wire [0:0] m_axi_gmem_2_WREADY,
	output wire [63:0] m_axi_gmem_2_WSTRB,
	output wire [0:0] m_axi_gmem_2_WVALID,
	output wire [63:0] m_axi_gmem_3_ARADDR,
	output wire [1:0] m_axi_gmem_3_ARBURST,
	output wire [3:0] m_axi_gmem_3_ARCACHE,
	output wire [0:0] m_axi_gmem_3_ARID,
	output wire [7:0] m_axi_gmem_3_ARLEN,
	output wire [1:0] m_axi_gmem_3_ARLOCK,
	output wire [2:0] m_axi_gmem_3_ARPROT,
	output wire [3:0] m_axi_gmem_3_ARQOS,
	input wire [0:0] m_axi_gmem_3_ARREADY,
	output wire [3:0] m_axi_gmem_3_ARREGION,
	output wire [2:0] m_axi_gmem_3_ARSIZE,
	output wire [0:0] m_axi_gmem_3_ARVALID,
	output wire [63:0] m_axi_gmem_3_AWADDR,
	output wire [1:0] m_axi_gmem_3_AWBURST,
	output wire [3:0] m_axi_gmem_3_AWCACHE,
	output wire [0:0] m_axi_gmem_3_AWID,
	output wire [7:0] m_axi_gmem_3_AWLEN,
	output wire [1:0] m_axi_gmem_3_AWLOCK,
	output wire [2:0] m_axi_gmem_3_AWPROT,
	output wire [3:0] m_axi_gmem_3_AWQOS,
	input wire [0:0] m_axi_gmem_3_AWREADY,
	output wire [3:0] m_axi_gmem_3_AWREGION,
	output wire [2:0] m_axi_gmem_3_AWSIZE,
	output wire [0:0] m_axi_gmem_3_AWVALID,
	input wire [0:0] m_axi_gmem_3_BID,
	output wire [0:0] m_axi_gmem_3_BREADY,
	input wire [1:0] m_axi_gmem_3_BRESP,
	input wire [0:0] m_axi_gmem_3_BVALID,
	input wire [511:0] m_axi_gmem_3_RDATA,
	input wire [0:0] m_axi_gmem_3_RID,
	input wire [0:0] m_axi_gmem_3_RLAST,
	output wire [0:0] m_axi_gmem_3_RREADY,
	input wire [1:0] m_axi_gmem_3_RRESP,
	input wire [0:0] m_axi_gmem_3_RVALID,
	output wire [511:0] m_axi_gmem_3_WDATA,
	output wire [0:0] m_axi_gmem_3_WLAST,
	input wire [0:0] m_axi_gmem_3_WREADY,
	output wire [63:0] m_axi_gmem_3_WSTRB,
	output wire [0:0] m_axi_gmem_3_WVALID,
	output wire [63:0] m_axi_gmem_4_ARADDR,
	output wire [1:0] m_axi_gmem_4_ARBURST,
	output wire [3:0] m_axi_gmem_4_ARCACHE,
	output wire [0:0] m_axi_gmem_4_ARID,
	output wire [7:0] m_axi_gmem_4_ARLEN,
	output wire [1:0] m_axi_gmem_4_ARLOCK,
	output wire [2:0] m_axi_gmem_4_ARPROT,
	output wire [3:0] m_axi_gmem_4_ARQOS,
	input wire [0:0] m_axi_gmem_4_ARREADY,
	output wire [3:0] m_axi_gmem_4_ARREGION,
	output wire [2:0] m_axi_gmem_4_ARSIZE,
	output wire [0:0] m_axi_gmem_4_ARVALID,
	output wire [63:0] m_axi_gmem_4_AWADDR,
	output wire [1:0] m_axi_gmem_4_AWBURST,
	output wire [3:0] m_axi_gmem_4_AWCACHE,
	output wire [0:0] m_axi_gmem_4_AWID,
	output wire [7:0] m_axi_gmem_4_AWLEN,
	output wire [1:0] m_axi_gmem_4_AWLOCK,
	output wire [2:0] m_axi_gmem_4_AWPROT,
	output wire [3:0] m_axi_gmem_4_AWQOS,
	input wire [0:0] m_axi_gmem_4_AWREADY,
	output wire [3:0] m_axi_gmem_4_AWREGION,
	output wire [2:0] m_axi_gmem_4_AWSIZE,
	output wire [0:0] m_axi_gmem_4_AWVALID,
	input wire [0:0] m_axi_gmem_4_BID,
	output wire [0:0] m_axi_gmem_4_BREADY,
	input wire [1:0] m_axi_gmem_4_BRESP,
	input wire [0:0] m_axi_gmem_4_BVALID,
	input wire [511:0] m_axi_gmem_4_RDATA,
	input wire [0:0] m_axi_gmem_4_RID,
	input wire [0:0] m_axi_gmem_4_RLAST,
	output wire [0:0] m_axi_gmem_4_RREADY,
	input wire [1:0] m_axi_gmem_4_RRESP,
	input wire [0:0] m_axi_gmem_4_RVALID,
	output wire [511:0] m_axi_gmem_4_WDATA,
	output wire [0:0] m_axi_gmem_4_WLAST,
	input wire [0:0] m_axi_gmem_4_WREADY,
	output wire [63:0] m_axi_gmem_4_WSTRB,
	output wire [0:0] m_axi_gmem_4_WVALID,
	output wire [63:0] m_axi_gmem_5_ARADDR,
	output wire [1:0] m_axi_gmem_5_ARBURST,
	output wire [3:0] m_axi_gmem_5_ARCACHE,
	output wire [0:0] m_axi_gmem_5_ARID,
	output wire [7:0] m_axi_gmem_5_ARLEN,
	output wire [1:0] m_axi_gmem_5_ARLOCK,
	output wire [2:0] m_axi_gmem_5_ARPROT,
	output wire [3:0] m_axi_gmem_5_ARQOS,
	input wire [0:0] m_axi_gmem_5_ARREADY,
	output wire [3:0] m_axi_gmem_5_ARREGION,
	output wire [2:0] m_axi_gmem_5_ARSIZE,
	output wire [0:0] m_axi_gmem_5_ARVALID,
	output wire [63:0] m_axi_gmem_5_AWADDR,
	output wire [1:0] m_axi_gmem_5_AWBURST,
	output wire [3:0] m_axi_gmem_5_AWCACHE,
	output wire [0:0] m_axi_gmem_5_AWID,
	output wire [7:0] m_axi_gmem_5_AWLEN,
	output wire [1:0] m_axi_gmem_5_AWLOCK,
	output wire [2:0] m_axi_gmem_5_AWPROT,
	output wire [3:0] m_axi_gmem_5_AWQOS,
	input wire [0:0] m_axi_gmem_5_AWREADY,
	output wire [3:0] m_axi_gmem_5_AWREGION,
	output wire [2:0] m_axi_gmem_5_AWSIZE,
	output wire [0:0] m_axi_gmem_5_AWVALID,
	input wire [0:0] m_axi_gmem_5_BID,
	output wire [0:0] m_axi_gmem_5_BREADY,
	input wire [1:0] m_axi_gmem_5_BRESP,
	input wire [0:0] m_axi_gmem_5_BVALID,
	input wire [511:0] m_axi_gmem_5_RDATA,
	input wire [0:0] m_axi_gmem_5_RID,
	input wire [0:0] m_axi_gmem_5_RLAST,
	output wire [0:0] m_axi_gmem_5_RREADY,
	input wire [1:0] m_axi_gmem_5_RRESP,
	input wire [0:0] m_axi_gmem_5_RVALID,
	output wire [511:0] m_axi_gmem_5_WDATA,
	output wire [0:0] m_axi_gmem_5_WLAST,
	input wire [0:0] m_axi_gmem_5_WREADY,
	output wire [63:0] m_axi_gmem_5_WSTRB,
	output wire [0:0] m_axi_gmem_5_WVALID,
	output wire [63:0] m_axi_gmem_6_ARADDR,
	output wire [1:0] m_axi_gmem_6_ARBURST,
	output wire [3:0] m_axi_gmem_6_ARCACHE,
	output wire [0:0] m_axi_gmem_6_ARID,
	output wire [7:0] m_axi_gmem_6_ARLEN,
	output wire [1:0] m_axi_gmem_6_ARLOCK,
	output wire [2:0] m_axi_gmem_6_ARPROT,
	output wire [3:0] m_axi_gmem_6_ARQOS,
	input wire [0:0] m_axi_gmem_6_ARREADY,
	output wire [3:0] m_axi_gmem_6_ARREGION,
	output wire [2:0] m_axi_gmem_6_ARSIZE,
	output wire [0:0] m_axi_gmem_6_ARVALID,
	output wire [63:0] m_axi_gmem_6_AWADDR,
	output wire [1:0] m_axi_gmem_6_AWBURST,
	output wire [3:0] m_axi_gmem_6_AWCACHE,
	output wire [0:0] m_axi_gmem_6_AWID,
	output wire [7:0] m_axi_gmem_6_AWLEN,
	output wire [1:0] m_axi_gmem_6_AWLOCK,
	output wire [2:0] m_axi_gmem_6_AWPROT,
	output wire [3:0] m_axi_gmem_6_AWQOS,
	input wire [0:0] m_axi_gmem_6_AWREADY,
	output wire [3:0] m_axi_gmem_6_AWREGION,
	output wire [2:0] m_axi_gmem_6_AWSIZE,
	output wire [0:0] m_axi_gmem_6_AWVALID,
	input wire [0:0] m_axi_gmem_6_BID,
	output wire [0:0] m_axi_gmem_6_BREADY,
	input wire [1:0] m_axi_gmem_6_BRESP,
	input wire [0:0] m_axi_gmem_6_BVALID,
	input wire [511:0] m_axi_gmem_6_RDATA,
	input wire [0:0] m_axi_gmem_6_RID,
	input wire [0:0] m_axi_gmem_6_RLAST,
	output wire [0:0] m_axi_gmem_6_RREADY,
	input wire [1:0] m_axi_gmem_6_RRESP,
	input wire [0:0] m_axi_gmem_6_RVALID,
	output wire [511:0] m_axi_gmem_6_WDATA,
	output wire [0:0] m_axi_gmem_6_WLAST,
	input wire [0:0] m_axi_gmem_6_WREADY,
	output wire [63:0] m_axi_gmem_6_WSTRB,
	output wire [0:0] m_axi_gmem_6_WVALID,
	output wire [63:0] m_axi_gmem_7_ARADDR,
	output wire [1:0] m_axi_gmem_7_ARBURST,
	output wire [3:0] m_axi_gmem_7_ARCACHE,
	output wire [0:0] m_axi_gmem_7_ARID,
	output wire [7:0] m_axi_gmem_7_ARLEN,
	output wire [1:0] m_axi_gmem_7_ARLOCK,
	output wire [2:0] m_axi_gmem_7_ARPROT,
	output wire [3:0] m_axi_gmem_7_ARQOS,
	input wire [0:0] m_axi_gmem_7_ARREADY,
	output wire [3:0] m_axi_gmem_7_ARREGION,
	output wire [2:0] m_axi_gmem_7_ARSIZE,
	output wire [0:0] m_axi_gmem_7_ARVALID,
	output wire [63:0] m_axi_gmem_7_AWADDR,
	output wire [1:0] m_axi_gmem_7_AWBURST,
	output wire [3:0] m_axi_gmem_7_AWCACHE,
	output wire [0:0] m_axi_gmem_7_AWID,
	output wire [7:0] m_axi_gmem_7_AWLEN,
	output wire [1:0] m_axi_gmem_7_AWLOCK,
	output wire [2:0] m_axi_gmem_7_AWPROT,
	output wire [3:0] m_axi_gmem_7_AWQOS,
	input wire [0:0] m_axi_gmem_7_AWREADY,
	output wire [3:0] m_axi_gmem_7_AWREGION,
	output wire [2:0] m_axi_gmem_7_AWSIZE,
	output wire [0:0] m_axi_gmem_7_AWVALID,
	input wire [0:0] m_axi_gmem_7_BID,
	output wire [0:0] m_axi_gmem_7_BREADY,
	input wire [1:0] m_axi_gmem_7_BRESP,
	input wire [0:0] m_axi_gmem_7_BVALID,
	input wire [511:0] m_axi_gmem_7_RDATA,
	input wire [0:0] m_axi_gmem_7_RID,
	input wire [0:0] m_axi_gmem_7_RLAST,
	output wire [0:0] m_axi_gmem_7_RREADY,
	input wire [1:0] m_axi_gmem_7_RRESP,
	input wire [0:0] m_axi_gmem_7_RVALID,
	output wire [511:0] m_axi_gmem_7_WDATA,
	output wire [0:0] m_axi_gmem_7_WLAST,
	input wire [0:0] m_axi_gmem_7_WREADY,
	output wire [63:0] m_axi_gmem_7_WSTRB,
	output wire [0:0] m_axi_gmem_7_WVALID,
	output wire [63:0] p0_TDATA,
	input wire [0:0] p0_TREADY,
	output wire [0:0] p0_TVALID,
	output wire [63:0] p1_TDATA,
	input wire [0:0] p1_TREADY,
	output wire [0:0] p1_TVALID,
	output wire [63:0] p2_TDATA,
	input wire [0:0] p2_TREADY,
	output wire [0:0] p2_TVALID,
	output wire [63:0] p3_TDATA,
	input wire [0:0] p3_TREADY,
	output wire [0:0] p3_TVALID,
	output wire [63:0] p4_TDATA,
	input wire [0:0] p4_TREADY,
	output wire [0:0] p4_TVALID,
	output wire [63:0] p5_TDATA,
	input wire [0:0] p5_TREADY,
	output wire [0:0] p5_TVALID,
	output wire [63:0] p6_TDATA,
	input wire [0:0] p6_TREADY,
	output wire [0:0] p6_TVALID,
	output wire [63:0] p7_TDATA,
	input wire [0:0] p7_TREADY,
	output wire [0:0] p7_TVALID,
	input wire [31:0] s_axi_control_ARADDR,
	output wire [0:0] s_axi_control_ARREADY,
	input wire [0:0] s_axi_control_ARVALID,
	input wire [31:0] s_axi_control_AWADDR,
	output wire [0:0] s_axi_control_AWREADY,
	input wire [0:0] s_axi_control_AWVALID,
	input wire [0:0] s_axi_control_BREADY,
	output wire [1:0] s_axi_control_BRESP,
	output wire [0:0] s_axi_control_BVALID,
	output wire [31:0] s_axi_control_RDATA,
	input wire [0:0] s_axi_control_RREADY,
	output wire [1:0] s_axi_control_RRESP,
	output wire [0:0] s_axi_control_RVALID,
	input wire [31:0] s_axi_control_WDATA,
	output wire [0:0] s_axi_control_WREADY,
	input wire [3:0] s_axi_control_WSTRB,
	input wire [0:0] s_axi_control_WVALID
);


krnl_hll_rtl_int krnl_hll_rtl_int_inst0 (
	.ap_aclk (ap_clk),
	.ap_aclk_2 (ap_clk_2),
	.ap_rst_n (ap_rst_n),
	.ap_rst_n_2 (ap_rst_n_2),
	.m_axi_gmem_0_ARADDR (m_axi_gmem_0_ARADDR),
	.m_axi_gmem_0_ARBURST (m_axi_gmem_0_ARBURST),
	.m_axi_gmem_0_ARCACHE (m_axi_gmem_0_ARCACHE),
	.m_axi_gmem_0_ARID (m_axi_gmem_0_ARID),
	.m_axi_gmem_0_ARLEN (m_axi_gmem_0_ARLEN),
	.m_axi_gmem_0_ARLOCK (m_axi_gmem_0_ARLOCK),
	.m_axi_gmem_0_ARPROT (m_axi_gmem_0_ARPROT),
	.m_axi_gmem_0_ARQOS (m_axi_gmem_0_ARQOS),
	.m_axi_gmem_0_ARREADY (m_axi_gmem_0_ARREADY),
	.m_axi_gmem_0_ARREGION (m_axi_gmem_0_ARREGION),
	.m_axi_gmem_0_ARSIZE (m_axi_gmem_0_ARSIZE),
	.m_axi_gmem_0_ARVALID (m_axi_gmem_0_ARVALID),
	.m_axi_gmem_0_AWADDR (m_axi_gmem_0_AWADDR),
	.m_axi_gmem_0_AWBURST (m_axi_gmem_0_AWBURST),
	.m_axi_gmem_0_AWCACHE (m_axi_gmem_0_AWCACHE),
	.m_axi_gmem_0_AWID (m_axi_gmem_0_AWID),
	.m_axi_gmem_0_AWLEN (m_axi_gmem_0_AWLEN),
	.m_axi_gmem_0_AWLOCK (m_axi_gmem_0_AWLOCK),
	.m_axi_gmem_0_AWPROT (m_axi_gmem_0_AWPROT),
	.m_axi_gmem_0_AWQOS (m_axi_gmem_0_AWQOS),
	.m_axi_gmem_0_AWREADY (m_axi_gmem_0_AWREADY),
	.m_axi_gmem_0_AWREGION (m_axi_gmem_0_AWREGION),
	.m_axi_gmem_0_AWSIZE (m_axi_gmem_0_AWSIZE),
	.m_axi_gmem_0_AWVALID (m_axi_gmem_0_AWVALID),
	.m_axi_gmem_0_BID (m_axi_gmem_0_BID),
	.m_axi_gmem_0_BREADY (m_axi_gmem_0_BREADY),
	.m_axi_gmem_0_BRESP (m_axi_gmem_0_BRESP),
	.m_axi_gmem_0_BVALID (m_axi_gmem_0_BVALID),
	.m_axi_gmem_0_RDATA (m_axi_gmem_0_RDATA),
	.m_axi_gmem_0_RID (m_axi_gmem_0_RID),
	.m_axi_gmem_0_RLAST (m_axi_gmem_0_RLAST),
	.m_axi_gmem_0_RREADY (m_axi_gmem_0_RREADY),
	.m_axi_gmem_0_RRESP (m_axi_gmem_0_RRESP),
	.m_axi_gmem_0_RVALID (m_axi_gmem_0_RVALID),
	.m_axi_gmem_0_WDATA (m_axi_gmem_0_WDATA),
	.m_axi_gmem_0_WLAST (m_axi_gmem_0_WLAST),
	.m_axi_gmem_0_WREADY (m_axi_gmem_0_WREADY),
	.m_axi_gmem_0_WSTRB (m_axi_gmem_0_WSTRB),
	.m_axi_gmem_0_WVALID (m_axi_gmem_0_WVALID),
	.m_axi_gmem_1_ARADDR (m_axi_gmem_1_ARADDR),
	.m_axi_gmem_1_ARBURST (m_axi_gmem_1_ARBURST),
	.m_axi_gmem_1_ARCACHE (m_axi_gmem_1_ARCACHE),
	.m_axi_gmem_1_ARID (m_axi_gmem_1_ARID),
	.m_axi_gmem_1_ARLEN (m_axi_gmem_1_ARLEN),
	.m_axi_gmem_1_ARLOCK (m_axi_gmem_1_ARLOCK),
	.m_axi_gmem_1_ARPROT (m_axi_gmem_1_ARPROT),
	.m_axi_gmem_1_ARQOS (m_axi_gmem_1_ARQOS),
	.m_axi_gmem_1_ARREADY (m_axi_gmem_1_ARREADY),
	.m_axi_gmem_1_ARREGION (m_axi_gmem_1_ARREGION),
	.m_axi_gmem_1_ARSIZE (m_axi_gmem_1_ARSIZE),
	.m_axi_gmem_1_ARVALID (m_axi_gmem_1_ARVALID),
	.m_axi_gmem_1_AWADDR (m_axi_gmem_1_AWADDR),
	.m_axi_gmem_1_AWBURST (m_axi_gmem_1_AWBURST),
	.m_axi_gmem_1_AWCACHE (m_axi_gmem_1_AWCACHE),
	.m_axi_gmem_1_AWID (m_axi_gmem_1_AWID),
	.m_axi_gmem_1_AWLEN (m_axi_gmem_1_AWLEN),
	.m_axi_gmem_1_AWLOCK (m_axi_gmem_1_AWLOCK),
	.m_axi_gmem_1_AWPROT (m_axi_gmem_1_AWPROT),
	.m_axi_gmem_1_AWQOS (m_axi_gmem_1_AWQOS),
	.m_axi_gmem_1_AWREADY (m_axi_gmem_1_AWREADY),
	.m_axi_gmem_1_AWREGION (m_axi_gmem_1_AWREGION),
	.m_axi_gmem_1_AWSIZE (m_axi_gmem_1_AWSIZE),
	.m_axi_gmem_1_AWVALID (m_axi_gmem_1_AWVALID),
	.m_axi_gmem_1_BID (m_axi_gmem_1_BID),
	.m_axi_gmem_1_BREADY (m_axi_gmem_1_BREADY),
	.m_axi_gmem_1_BRESP (m_axi_gmem_1_BRESP),
	.m_axi_gmem_1_BVALID (m_axi_gmem_1_BVALID),
	.m_axi_gmem_1_RDATA (m_axi_gmem_1_RDATA),
	.m_axi_gmem_1_RID (m_axi_gmem_1_RID),
	.m_axi_gmem_1_RLAST (m_axi_gmem_1_RLAST),
	.m_axi_gmem_1_RREADY (m_axi_gmem_1_RREADY),
	.m_axi_gmem_1_RRESP (m_axi_gmem_1_RRESP),
	.m_axi_gmem_1_RVALID (m_axi_gmem_1_RVALID),
	.m_axi_gmem_1_WDATA (m_axi_gmem_1_WDATA),
	.m_axi_gmem_1_WLAST (m_axi_gmem_1_WLAST),
	.m_axi_gmem_1_WREADY (m_axi_gmem_1_WREADY),
	.m_axi_gmem_1_WSTRB (m_axi_gmem_1_WSTRB),
	.m_axi_gmem_1_WVALID (m_axi_gmem_1_WVALID),
	.m_axi_gmem_2_ARADDR (m_axi_gmem_2_ARADDR),
	.m_axi_gmem_2_ARBURST (m_axi_gmem_2_ARBURST),
	.m_axi_gmem_2_ARCACHE (m_axi_gmem_2_ARCACHE),
	.m_axi_gmem_2_ARID (m_axi_gmem_2_ARID),
	.m_axi_gmem_2_ARLEN (m_axi_gmem_2_ARLEN),
	.m_axi_gmem_2_ARLOCK (m_axi_gmem_2_ARLOCK),
	.m_axi_gmem_2_ARPROT (m_axi_gmem_2_ARPROT),
	.m_axi_gmem_2_ARQOS (m_axi_gmem_2_ARQOS),
	.m_axi_gmem_2_ARREADY (m_axi_gmem_2_ARREADY),
	.m_axi_gmem_2_ARREGION (m_axi_gmem_2_ARREGION),
	.m_axi_gmem_2_ARSIZE (m_axi_gmem_2_ARSIZE),
	.m_axi_gmem_2_ARVALID (m_axi_gmem_2_ARVALID),
	.m_axi_gmem_2_AWADDR (m_axi_gmem_2_AWADDR),
	.m_axi_gmem_2_AWBURST (m_axi_gmem_2_AWBURST),
	.m_axi_gmem_2_AWCACHE (m_axi_gmem_2_AWCACHE),
	.m_axi_gmem_2_AWID (m_axi_gmem_2_AWID),
	.m_axi_gmem_2_AWLEN (m_axi_gmem_2_AWLEN),
	.m_axi_gmem_2_AWLOCK (m_axi_gmem_2_AWLOCK),
	.m_axi_gmem_2_AWPROT (m_axi_gmem_2_AWPROT),
	.m_axi_gmem_2_AWQOS (m_axi_gmem_2_AWQOS),
	.m_axi_gmem_2_AWREADY (m_axi_gmem_2_AWREADY),
	.m_axi_gmem_2_AWREGION (m_axi_gmem_2_AWREGION),
	.m_axi_gmem_2_AWSIZE (m_axi_gmem_2_AWSIZE),
	.m_axi_gmem_2_AWVALID (m_axi_gmem_2_AWVALID),
	.m_axi_gmem_2_BID (m_axi_gmem_2_BID),
	.m_axi_gmem_2_BREADY (m_axi_gmem_2_BREADY),
	.m_axi_gmem_2_BRESP (m_axi_gmem_2_BRESP),
	.m_axi_gmem_2_BVALID (m_axi_gmem_2_BVALID),
	.m_axi_gmem_2_RDATA (m_axi_gmem_2_RDATA),
	.m_axi_gmem_2_RID (m_axi_gmem_2_RID),
	.m_axi_gmem_2_RLAST (m_axi_gmem_2_RLAST),
	.m_axi_gmem_2_RREADY (m_axi_gmem_2_RREADY),
	.m_axi_gmem_2_RRESP (m_axi_gmem_2_RRESP),
	.m_axi_gmem_2_RVALID (m_axi_gmem_2_RVALID),
	.m_axi_gmem_2_WDATA (m_axi_gmem_2_WDATA),
	.m_axi_gmem_2_WLAST (m_axi_gmem_2_WLAST),
	.m_axi_gmem_2_WREADY (m_axi_gmem_2_WREADY),
	.m_axi_gmem_2_WSTRB (m_axi_gmem_2_WSTRB),
	.m_axi_gmem_2_WVALID (m_axi_gmem_2_WVALID),
	.m_axi_gmem_3_ARADDR (m_axi_gmem_3_ARADDR),
	.m_axi_gmem_3_ARBURST (m_axi_gmem_3_ARBURST),
	.m_axi_gmem_3_ARCACHE (m_axi_gmem_3_ARCACHE),
	.m_axi_gmem_3_ARID (m_axi_gmem_3_ARID),
	.m_axi_gmem_3_ARLEN (m_axi_gmem_3_ARLEN),
	.m_axi_gmem_3_ARLOCK (m_axi_gmem_3_ARLOCK),
	.m_axi_gmem_3_ARPROT (m_axi_gmem_3_ARPROT),
	.m_axi_gmem_3_ARQOS (m_axi_gmem_3_ARQOS),
	.m_axi_gmem_3_ARREADY (m_axi_gmem_3_ARREADY),
	.m_axi_gmem_3_ARREGION (m_axi_gmem_3_ARREGION),
	.m_axi_gmem_3_ARSIZE (m_axi_gmem_3_ARSIZE),
	.m_axi_gmem_3_ARVALID (m_axi_gmem_3_ARVALID),
	.m_axi_gmem_3_AWADDR (m_axi_gmem_3_AWADDR),
	.m_axi_gmem_3_AWBURST (m_axi_gmem_3_AWBURST),
	.m_axi_gmem_3_AWCACHE (m_axi_gmem_3_AWCACHE),
	.m_axi_gmem_3_AWID (m_axi_gmem_3_AWID),
	.m_axi_gmem_3_AWLEN (m_axi_gmem_3_AWLEN),
	.m_axi_gmem_3_AWLOCK (m_axi_gmem_3_AWLOCK),
	.m_axi_gmem_3_AWPROT (m_axi_gmem_3_AWPROT),
	.m_axi_gmem_3_AWQOS (m_axi_gmem_3_AWQOS),
	.m_axi_gmem_3_AWREADY (m_axi_gmem_3_AWREADY),
	.m_axi_gmem_3_AWREGION (m_axi_gmem_3_AWREGION),
	.m_axi_gmem_3_AWSIZE (m_axi_gmem_3_AWSIZE),
	.m_axi_gmem_3_AWVALID (m_axi_gmem_3_AWVALID),
	.m_axi_gmem_3_BID (m_axi_gmem_3_BID),
	.m_axi_gmem_3_BREADY (m_axi_gmem_3_BREADY),
	.m_axi_gmem_3_BRESP (m_axi_gmem_3_BRESP),
	.m_axi_gmem_3_BVALID (m_axi_gmem_3_BVALID),
	.m_axi_gmem_3_RDATA (m_axi_gmem_3_RDATA),
	.m_axi_gmem_3_RID (m_axi_gmem_3_RID),
	.m_axi_gmem_3_RLAST (m_axi_gmem_3_RLAST),
	.m_axi_gmem_3_RREADY (m_axi_gmem_3_RREADY),
	.m_axi_gmem_3_RRESP (m_axi_gmem_3_RRESP),
	.m_axi_gmem_3_RVALID (m_axi_gmem_3_RVALID),
	.m_axi_gmem_3_WDATA (m_axi_gmem_3_WDATA),
	.m_axi_gmem_3_WLAST (m_axi_gmem_3_WLAST),
	.m_axi_gmem_3_WREADY (m_axi_gmem_3_WREADY),
	.m_axi_gmem_3_WSTRB (m_axi_gmem_3_WSTRB),
	.m_axi_gmem_3_WVALID (m_axi_gmem_3_WVALID),
	.m_axi_gmem_4_ARADDR (m_axi_gmem_4_ARADDR),
	.m_axi_gmem_4_ARBURST (m_axi_gmem_4_ARBURST),
	.m_axi_gmem_4_ARCACHE (m_axi_gmem_4_ARCACHE),
	.m_axi_gmem_4_ARID (m_axi_gmem_4_ARID),
	.m_axi_gmem_4_ARLEN (m_axi_gmem_4_ARLEN),
	.m_axi_gmem_4_ARLOCK (m_axi_gmem_4_ARLOCK),
	.m_axi_gmem_4_ARPROT (m_axi_gmem_4_ARPROT),
	.m_axi_gmem_4_ARQOS (m_axi_gmem_4_ARQOS),
	.m_axi_gmem_4_ARREADY (m_axi_gmem_4_ARREADY),
	.m_axi_gmem_4_ARREGION (m_axi_gmem_4_ARREGION),
	.m_axi_gmem_4_ARSIZE (m_axi_gmem_4_ARSIZE),
	.m_axi_gmem_4_ARVALID (m_axi_gmem_4_ARVALID),
	.m_axi_gmem_4_AWADDR (m_axi_gmem_4_AWADDR),
	.m_axi_gmem_4_AWBURST (m_axi_gmem_4_AWBURST),
	.m_axi_gmem_4_AWCACHE (m_axi_gmem_4_AWCACHE),
	.m_axi_gmem_4_AWID (m_axi_gmem_4_AWID),
	.m_axi_gmem_4_AWLEN (m_axi_gmem_4_AWLEN),
	.m_axi_gmem_4_AWLOCK (m_axi_gmem_4_AWLOCK),
	.m_axi_gmem_4_AWPROT (m_axi_gmem_4_AWPROT),
	.m_axi_gmem_4_AWQOS (m_axi_gmem_4_AWQOS),
	.m_axi_gmem_4_AWREADY (m_axi_gmem_4_AWREADY),
	.m_axi_gmem_4_AWREGION (m_axi_gmem_4_AWREGION),
	.m_axi_gmem_4_AWSIZE (m_axi_gmem_4_AWSIZE),
	.m_axi_gmem_4_AWVALID (m_axi_gmem_4_AWVALID),
	.m_axi_gmem_4_BID (m_axi_gmem_4_BID),
	.m_axi_gmem_4_BREADY (m_axi_gmem_4_BREADY),
	.m_axi_gmem_4_BRESP (m_axi_gmem_4_BRESP),
	.m_axi_gmem_4_BVALID (m_axi_gmem_4_BVALID),
	.m_axi_gmem_4_RDATA (m_axi_gmem_4_RDATA),
	.m_axi_gmem_4_RID (m_axi_gmem_4_RID),
	.m_axi_gmem_4_RLAST (m_axi_gmem_4_RLAST),
	.m_axi_gmem_4_RREADY (m_axi_gmem_4_RREADY),
	.m_axi_gmem_4_RRESP (m_axi_gmem_4_RRESP),
	.m_axi_gmem_4_RVALID (m_axi_gmem_4_RVALID),
	.m_axi_gmem_4_WDATA (m_axi_gmem_4_WDATA),
	.m_axi_gmem_4_WLAST (m_axi_gmem_4_WLAST),
	.m_axi_gmem_4_WREADY (m_axi_gmem_4_WREADY),
	.m_axi_gmem_4_WSTRB (m_axi_gmem_4_WSTRB),
	.m_axi_gmem_4_WVALID (m_axi_gmem_4_WVALID),
	.m_axi_gmem_5_ARADDR (m_axi_gmem_5_ARADDR),
	.m_axi_gmem_5_ARBURST (m_axi_gmem_5_ARBURST),
	.m_axi_gmem_5_ARCACHE (m_axi_gmem_5_ARCACHE),
	.m_axi_gmem_5_ARID (m_axi_gmem_5_ARID),
	.m_axi_gmem_5_ARLEN (m_axi_gmem_5_ARLEN),
	.m_axi_gmem_5_ARLOCK (m_axi_gmem_5_ARLOCK),
	.m_axi_gmem_5_ARPROT (m_axi_gmem_5_ARPROT),
	.m_axi_gmem_5_ARQOS (m_axi_gmem_5_ARQOS),
	.m_axi_gmem_5_ARREADY (m_axi_gmem_5_ARREADY),
	.m_axi_gmem_5_ARREGION (m_axi_gmem_5_ARREGION),
	.m_axi_gmem_5_ARSIZE (m_axi_gmem_5_ARSIZE),
	.m_axi_gmem_5_ARVALID (m_axi_gmem_5_ARVALID),
	.m_axi_gmem_5_AWADDR (m_axi_gmem_5_AWADDR),
	.m_axi_gmem_5_AWBURST (m_axi_gmem_5_AWBURST),
	.m_axi_gmem_5_AWCACHE (m_axi_gmem_5_AWCACHE),
	.m_axi_gmem_5_AWID (m_axi_gmem_5_AWID),
	.m_axi_gmem_5_AWLEN (m_axi_gmem_5_AWLEN),
	.m_axi_gmem_5_AWLOCK (m_axi_gmem_5_AWLOCK),
	.m_axi_gmem_5_AWPROT (m_axi_gmem_5_AWPROT),
	.m_axi_gmem_5_AWQOS (m_axi_gmem_5_AWQOS),
	.m_axi_gmem_5_AWREADY (m_axi_gmem_5_AWREADY),
	.m_axi_gmem_5_AWREGION (m_axi_gmem_5_AWREGION),
	.m_axi_gmem_5_AWSIZE (m_axi_gmem_5_AWSIZE),
	.m_axi_gmem_5_AWVALID (m_axi_gmem_5_AWVALID),
	.m_axi_gmem_5_BID (m_axi_gmem_5_BID),
	.m_axi_gmem_5_BREADY (m_axi_gmem_5_BREADY),
	.m_axi_gmem_5_BRESP (m_axi_gmem_5_BRESP),
	.m_axi_gmem_5_BVALID (m_axi_gmem_5_BVALID),
	.m_axi_gmem_5_RDATA (m_axi_gmem_5_RDATA),
	.m_axi_gmem_5_RID (m_axi_gmem_5_RID),
	.m_axi_gmem_5_RLAST (m_axi_gmem_5_RLAST),
	.m_axi_gmem_5_RREADY (m_axi_gmem_5_RREADY),
	.m_axi_gmem_5_RRESP (m_axi_gmem_5_RRESP),
	.m_axi_gmem_5_RVALID (m_axi_gmem_5_RVALID),
	.m_axi_gmem_5_WDATA (m_axi_gmem_5_WDATA),
	.m_axi_gmem_5_WLAST (m_axi_gmem_5_WLAST),
	.m_axi_gmem_5_WREADY (m_axi_gmem_5_WREADY),
	.m_axi_gmem_5_WSTRB (m_axi_gmem_5_WSTRB),
	.m_axi_gmem_5_WVALID (m_axi_gmem_5_WVALID),
	.m_axi_gmem_6_ARADDR (m_axi_gmem_6_ARADDR),
	.m_axi_gmem_6_ARBURST (m_axi_gmem_6_ARBURST),
	.m_axi_gmem_6_ARCACHE (m_axi_gmem_6_ARCACHE),
	.m_axi_gmem_6_ARID (m_axi_gmem_6_ARID),
	.m_axi_gmem_6_ARLEN (m_axi_gmem_6_ARLEN),
	.m_axi_gmem_6_ARLOCK (m_axi_gmem_6_ARLOCK),
	.m_axi_gmem_6_ARPROT (m_axi_gmem_6_ARPROT),
	.m_axi_gmem_6_ARQOS (m_axi_gmem_6_ARQOS),
	.m_axi_gmem_6_ARREADY (m_axi_gmem_6_ARREADY),
	.m_axi_gmem_6_ARREGION (m_axi_gmem_6_ARREGION),
	.m_axi_gmem_6_ARSIZE (m_axi_gmem_6_ARSIZE),
	.m_axi_gmem_6_ARVALID (m_axi_gmem_6_ARVALID),
	.m_axi_gmem_6_AWADDR (m_axi_gmem_6_AWADDR),
	.m_axi_gmem_6_AWBURST (m_axi_gmem_6_AWBURST),
	.m_axi_gmem_6_AWCACHE (m_axi_gmem_6_AWCACHE),
	.m_axi_gmem_6_AWID (m_axi_gmem_6_AWID),
	.m_axi_gmem_6_AWLEN (m_axi_gmem_6_AWLEN),
	.m_axi_gmem_6_AWLOCK (m_axi_gmem_6_AWLOCK),
	.m_axi_gmem_6_AWPROT (m_axi_gmem_6_AWPROT),
	.m_axi_gmem_6_AWQOS (m_axi_gmem_6_AWQOS),
	.m_axi_gmem_6_AWREADY (m_axi_gmem_6_AWREADY),
	.m_axi_gmem_6_AWREGION (m_axi_gmem_6_AWREGION),
	.m_axi_gmem_6_AWSIZE (m_axi_gmem_6_AWSIZE),
	.m_axi_gmem_6_AWVALID (m_axi_gmem_6_AWVALID),
	.m_axi_gmem_6_BID (m_axi_gmem_6_BID),
	.m_axi_gmem_6_BREADY (m_axi_gmem_6_BREADY),
	.m_axi_gmem_6_BRESP (m_axi_gmem_6_BRESP),
	.m_axi_gmem_6_BVALID (m_axi_gmem_6_BVALID),
	.m_axi_gmem_6_RDATA (m_axi_gmem_6_RDATA),
	.m_axi_gmem_6_RID (m_axi_gmem_6_RID),
	.m_axi_gmem_6_RLAST (m_axi_gmem_6_RLAST),
	.m_axi_gmem_6_RREADY (m_axi_gmem_6_RREADY),
	.m_axi_gmem_6_RRESP (m_axi_gmem_6_RRESP),
	.m_axi_gmem_6_RVALID (m_axi_gmem_6_RVALID),
	.m_axi_gmem_6_WDATA (m_axi_gmem_6_WDATA),
	.m_axi_gmem_6_WLAST (m_axi_gmem_6_WLAST),
	.m_axi_gmem_6_WREADY (m_axi_gmem_6_WREADY),
	.m_axi_gmem_6_WSTRB (m_axi_gmem_6_WSTRB),
	.m_axi_gmem_6_WVALID (m_axi_gmem_6_WVALID),
	.m_axi_gmem_7_ARADDR (m_axi_gmem_7_ARADDR),
	.m_axi_gmem_7_ARBURST (m_axi_gmem_7_ARBURST),
	.m_axi_gmem_7_ARCACHE (m_axi_gmem_7_ARCACHE),
	.m_axi_gmem_7_ARID (m_axi_gmem_7_ARID),
	.m_axi_gmem_7_ARLEN (m_axi_gmem_7_ARLEN),
	.m_axi_gmem_7_ARLOCK (m_axi_gmem_7_ARLOCK),
	.m_axi_gmem_7_ARPROT (m_axi_gmem_7_ARPROT),
	.m_axi_gmem_7_ARQOS (m_axi_gmem_7_ARQOS),
	.m_axi_gmem_7_ARREADY (m_axi_gmem_7_ARREADY),
	.m_axi_gmem_7_ARREGION (m_axi_gmem_7_ARREGION),
	.m_axi_gmem_7_ARSIZE (m_axi_gmem_7_ARSIZE),
	.m_axi_gmem_7_ARVALID (m_axi_gmem_7_ARVALID),
	.m_axi_gmem_7_AWADDR (m_axi_gmem_7_AWADDR),
	.m_axi_gmem_7_AWBURST (m_axi_gmem_7_AWBURST),
	.m_axi_gmem_7_AWCACHE (m_axi_gmem_7_AWCACHE),
	.m_axi_gmem_7_AWID (m_axi_gmem_7_AWID),
	.m_axi_gmem_7_AWLEN (m_axi_gmem_7_AWLEN),
	.m_axi_gmem_7_AWLOCK (m_axi_gmem_7_AWLOCK),
	.m_axi_gmem_7_AWPROT (m_axi_gmem_7_AWPROT),
	.m_axi_gmem_7_AWQOS (m_axi_gmem_7_AWQOS),
	.m_axi_gmem_7_AWREADY (m_axi_gmem_7_AWREADY),
	.m_axi_gmem_7_AWREGION (m_axi_gmem_7_AWREGION),
	.m_axi_gmem_7_AWSIZE (m_axi_gmem_7_AWSIZE),
	.m_axi_gmem_7_AWVALID (m_axi_gmem_7_AWVALID),
	.m_axi_gmem_7_BID (m_axi_gmem_7_BID),
	.m_axi_gmem_7_BREADY (m_axi_gmem_7_BREADY),
	.m_axi_gmem_7_BRESP (m_axi_gmem_7_BRESP),
	.m_axi_gmem_7_BVALID (m_axi_gmem_7_BVALID),
	.m_axi_gmem_7_RDATA (m_axi_gmem_7_RDATA),
	.m_axi_gmem_7_RID (m_axi_gmem_7_RID),
	.m_axi_gmem_7_RLAST (m_axi_gmem_7_RLAST),
	.m_axi_gmem_7_RREADY (m_axi_gmem_7_RREADY),
	.m_axi_gmem_7_RRESP (m_axi_gmem_7_RRESP),
	.m_axi_gmem_7_RVALID (m_axi_gmem_7_RVALID),
	.m_axi_gmem_7_WDATA (m_axi_gmem_7_WDATA),
	.m_axi_gmem_7_WLAST (m_axi_gmem_7_WLAST),
	.m_axi_gmem_7_WREADY (m_axi_gmem_7_WREADY),
	.m_axi_gmem_7_WSTRB (m_axi_gmem_7_WSTRB),
	.m_axi_gmem_7_WVALID (m_axi_gmem_7_WVALID),
	.p0_TDATA (p0_TDATA),
	.p0_TREADY (p0_TREADY),
	.p0_TVALID (p0_TVALID),
	.p1_TDATA (p1_TDATA),
	.p1_TREADY (p1_TREADY),
	.p1_TVALID (p1_TVALID),
	.p2_TDATA (p2_TDATA),
	.p2_TREADY (p2_TREADY),
	.p2_TVALID (p2_TVALID),
	.p3_TDATA (p3_TDATA),
	.p3_TREADY (p3_TREADY),
	.p3_TVALID (p3_TVALID),
	.p4_TDATA (p4_TDATA),
	.p4_TREADY (p4_TREADY),
	.p4_TVALID (p4_TVALID),
	.p5_TDATA (p5_TDATA),
	.p5_TREADY (p5_TREADY),
	.p5_TVALID (p5_TVALID),
	.p6_TDATA (p6_TDATA),
	.p6_TREADY (p6_TREADY),
	.p6_TVALID (p6_TVALID),
	.p7_TDATA (p7_TDATA),
	.p7_TREADY (p7_TREADY),
	.p7_TVALID (p7_TVALID),
	.s_axi_control_ARADDR (s_axi_control_ARADDR),
	.s_axi_control_ARREADY (s_axi_control_ARREADY),
	.s_axi_control_ARVALID (s_axi_control_ARVALID),
	.s_axi_control_AWADDR (s_axi_control_AWADDR),
	.s_axi_control_AWREADY (s_axi_control_AWREADY),
	.s_axi_control_AWVALID (s_axi_control_AWVALID),
	.s_axi_control_BREADY (s_axi_control_BREADY),
	.s_axi_control_BRESP (s_axi_control_BRESP),
	.s_axi_control_BVALID (s_axi_control_BVALID),
	.s_axi_control_RDATA (s_axi_control_RDATA),
	.s_axi_control_RREADY (s_axi_control_RREADY),
	.s_axi_control_RRESP (s_axi_control_RRESP),
	.s_axi_control_RVALID (s_axi_control_RVALID),
	.s_axi_control_WDATA (s_axi_control_WDATA),
	.s_axi_control_WREADY (s_axi_control_WREADY),
	.s_axi_control_WSTRB (s_axi_control_WSTRB),
	.s_axi_control_WVALID (s_axi_control_WVALID)
);

endmodule

