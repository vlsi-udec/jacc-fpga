`timescale 1ns / 1ps

module hll_mem (
	output logic [0:0] busy_out,
	input logic [0:0] clk,
	input logic [3:0] data_0,
	input logic [3:0] data_1,
	input logic [3:0] data_2,
	input logic [3:0] data_3,
	input logic [3:0] data_4,
	input logic [3:0] data_5,
	input logic [3:0] data_6,
	input logic [3:0] data_7,
	input logic [13:0] idx_0,
	input logic [13:0] idx_1,
	input logic [13:0] idx_2,
	input logic [13:0] idx_3,
	input logic [13:0] idx_4,
	input logic [13:0] idx_5,
	input logic [13:0] idx_6,
	input logic [13:0] idx_7,
	input logic [0:0] last,
	output logic [511:0] out_data,
	input logic [0:0] out_ready,
	output logic [0:0] out_valid,
	input logic [7:0] valid
);

logic [63:0] out_mem[7:0];
logic [63:0] in_mem[7:0];
logic [9:0] r_idx[7:0];
logic [63:0] r_data[7:0];
logic [9:0] r2_idx[7:0];
logic [9:0] r3_idx[7:0];
logic [63:0] r2_data[7:0];
logic [63:0] r3_data[7:0];
logic [7:0] r_valid[2:0];
logic [9:0] mem_wr_addr[7:0];
logic [9:0] mem_rd_addr[7:0];
logic [63:0] max_tree_0[3:0];
logic [63:0] max_tree_1[1:0];
logic [63:0] max_tree_2[0:0];
logic [63:0] mem_0[1023:0];
logic [63:0] mem_1[1023:0];
logic [63:0] mem_2[1023:0];
logic [63:0] mem_3[1023:0];
logic [63:0] mem_4[1023:0];
logic [63:0] mem_5[1023:0];
logic [63:0] mem_6[1023:0];
logic [63:0] mem_7[1023:0];
logic [2:0] r_last = 3'd0;
logic [0:0] busy = 1'd0;
logic [9:0] out_cnt = 10'd0;
logic [3:0] out_mem_valid = 4'd0;
logic [0:0] reading_memory = 1'd0;
logic [0:0] out_valid_in;
logic [63:0] out_data_in;
logic [3:0] out_valid_cnt = 4'd0;

initial begin
	mem_0[0] = 64'd0;
	mem_0[1] = 64'd0;
	mem_0[2] = 64'd0;
	mem_0[3] = 64'd0;
	mem_0[4] = 64'd0;
	mem_0[5] = 64'd0;
	mem_0[6] = 64'd0;
	mem_0[7] = 64'd0;
	mem_0[8] = 64'd0;
	mem_0[9] = 64'd0;
	mem_0[10] = 64'd0;
	mem_0[11] = 64'd0;
	mem_0[12] = 64'd0;
	mem_0[13] = 64'd0;
	mem_0[14] = 64'd0;
	mem_0[15] = 64'd0;
	mem_0[16] = 64'd0;
	mem_0[17] = 64'd0;
	mem_0[18] = 64'd0;
	mem_0[19] = 64'd0;
	mem_0[20] = 64'd0;
	mem_0[21] = 64'd0;
	mem_0[22] = 64'd0;
	mem_0[23] = 64'd0;
	mem_0[24] = 64'd0;
	mem_0[25] = 64'd0;
	mem_0[26] = 64'd0;
	mem_0[27] = 64'd0;
	mem_0[28] = 64'd0;
	mem_0[29] = 64'd0;
	mem_0[30] = 64'd0;
	mem_0[31] = 64'd0;
	mem_0[32] = 64'd0;
	mem_0[33] = 64'd0;
	mem_0[34] = 64'd0;
	mem_0[35] = 64'd0;
	mem_0[36] = 64'd0;
	mem_0[37] = 64'd0;
	mem_0[38] = 64'd0;
	mem_0[39] = 64'd0;
	mem_0[40] = 64'd0;
	mem_0[41] = 64'd0;
	mem_0[42] = 64'd0;
	mem_0[43] = 64'd0;
	mem_0[44] = 64'd0;
	mem_0[45] = 64'd0;
	mem_0[46] = 64'd0;
	mem_0[47] = 64'd0;
	mem_0[48] = 64'd0;
	mem_0[49] = 64'd0;
	mem_0[50] = 64'd0;
	mem_0[51] = 64'd0;
	mem_0[52] = 64'd0;
	mem_0[53] = 64'd0;
	mem_0[54] = 64'd0;
	mem_0[55] = 64'd0;
	mem_0[56] = 64'd0;
	mem_0[57] = 64'd0;
	mem_0[58] = 64'd0;
	mem_0[59] = 64'd0;
	mem_0[60] = 64'd0;
	mem_0[61] = 64'd0;
	mem_0[62] = 64'd0;
	mem_0[63] = 64'd0;
	mem_0[64] = 64'd0;
	mem_0[65] = 64'd0;
	mem_0[66] = 64'd0;
	mem_0[67] = 64'd0;
	mem_0[68] = 64'd0;
	mem_0[69] = 64'd0;
	mem_0[70] = 64'd0;
	mem_0[71] = 64'd0;
	mem_0[72] = 64'd0;
	mem_0[73] = 64'd0;
	mem_0[74] = 64'd0;
	mem_0[75] = 64'd0;
	mem_0[76] = 64'd0;
	mem_0[77] = 64'd0;
	mem_0[78] = 64'd0;
	mem_0[79] = 64'd0;
	mem_0[80] = 64'd0;
	mem_0[81] = 64'd0;
	mem_0[82] = 64'd0;
	mem_0[83] = 64'd0;
	mem_0[84] = 64'd0;
	mem_0[85] = 64'd0;
	mem_0[86] = 64'd0;
	mem_0[87] = 64'd0;
	mem_0[88] = 64'd0;
	mem_0[89] = 64'd0;
	mem_0[90] = 64'd0;
	mem_0[91] = 64'd0;
	mem_0[92] = 64'd0;
	mem_0[93] = 64'd0;
	mem_0[94] = 64'd0;
	mem_0[95] = 64'd0;
	mem_0[96] = 64'd0;
	mem_0[97] = 64'd0;
	mem_0[98] = 64'd0;
	mem_0[99] = 64'd0;
	mem_0[100] = 64'd0;
	mem_0[101] = 64'd0;
	mem_0[102] = 64'd0;
	mem_0[103] = 64'd0;
	mem_0[104] = 64'd0;
	mem_0[105] = 64'd0;
	mem_0[106] = 64'd0;
	mem_0[107] = 64'd0;
	mem_0[108] = 64'd0;
	mem_0[109] = 64'd0;
	mem_0[110] = 64'd0;
	mem_0[111] = 64'd0;
	mem_0[112] = 64'd0;
	mem_0[113] = 64'd0;
	mem_0[114] = 64'd0;
	mem_0[115] = 64'd0;
	mem_0[116] = 64'd0;
	mem_0[117] = 64'd0;
	mem_0[118] = 64'd0;
	mem_0[119] = 64'd0;
	mem_0[120] = 64'd0;
	mem_0[121] = 64'd0;
	mem_0[122] = 64'd0;
	mem_0[123] = 64'd0;
	mem_0[124] = 64'd0;
	mem_0[125] = 64'd0;
	mem_0[126] = 64'd0;
	mem_0[127] = 64'd0;
	mem_0[128] = 64'd0;
	mem_0[129] = 64'd0;
	mem_0[130] = 64'd0;
	mem_0[131] = 64'd0;
	mem_0[132] = 64'd0;
	mem_0[133] = 64'd0;
	mem_0[134] = 64'd0;
	mem_0[135] = 64'd0;
	mem_0[136] = 64'd0;
	mem_0[137] = 64'd0;
	mem_0[138] = 64'd0;
	mem_0[139] = 64'd0;
	mem_0[140] = 64'd0;
	mem_0[141] = 64'd0;
	mem_0[142] = 64'd0;
	mem_0[143] = 64'd0;
	mem_0[144] = 64'd0;
	mem_0[145] = 64'd0;
	mem_0[146] = 64'd0;
	mem_0[147] = 64'd0;
	mem_0[148] = 64'd0;
	mem_0[149] = 64'd0;
	mem_0[150] = 64'd0;
	mem_0[151] = 64'd0;
	mem_0[152] = 64'd0;
	mem_0[153] = 64'd0;
	mem_0[154] = 64'd0;
	mem_0[155] = 64'd0;
	mem_0[156] = 64'd0;
	mem_0[157] = 64'd0;
	mem_0[158] = 64'd0;
	mem_0[159] = 64'd0;
	mem_0[160] = 64'd0;
	mem_0[161] = 64'd0;
	mem_0[162] = 64'd0;
	mem_0[163] = 64'd0;
	mem_0[164] = 64'd0;
	mem_0[165] = 64'd0;
	mem_0[166] = 64'd0;
	mem_0[167] = 64'd0;
	mem_0[168] = 64'd0;
	mem_0[169] = 64'd0;
	mem_0[170] = 64'd0;
	mem_0[171] = 64'd0;
	mem_0[172] = 64'd0;
	mem_0[173] = 64'd0;
	mem_0[174] = 64'd0;
	mem_0[175] = 64'd0;
	mem_0[176] = 64'd0;
	mem_0[177] = 64'd0;
	mem_0[178] = 64'd0;
	mem_0[179] = 64'd0;
	mem_0[180] = 64'd0;
	mem_0[181] = 64'd0;
	mem_0[182] = 64'd0;
	mem_0[183] = 64'd0;
	mem_0[184] = 64'd0;
	mem_0[185] = 64'd0;
	mem_0[186] = 64'd0;
	mem_0[187] = 64'd0;
	mem_0[188] = 64'd0;
	mem_0[189] = 64'd0;
	mem_0[190] = 64'd0;
	mem_0[191] = 64'd0;
	mem_0[192] = 64'd0;
	mem_0[193] = 64'd0;
	mem_0[194] = 64'd0;
	mem_0[195] = 64'd0;
	mem_0[196] = 64'd0;
	mem_0[197] = 64'd0;
	mem_0[198] = 64'd0;
	mem_0[199] = 64'd0;
	mem_0[200] = 64'd0;
	mem_0[201] = 64'd0;
	mem_0[202] = 64'd0;
	mem_0[203] = 64'd0;
	mem_0[204] = 64'd0;
	mem_0[205] = 64'd0;
	mem_0[206] = 64'd0;
	mem_0[207] = 64'd0;
	mem_0[208] = 64'd0;
	mem_0[209] = 64'd0;
	mem_0[210] = 64'd0;
	mem_0[211] = 64'd0;
	mem_0[212] = 64'd0;
	mem_0[213] = 64'd0;
	mem_0[214] = 64'd0;
	mem_0[215] = 64'd0;
	mem_0[216] = 64'd0;
	mem_0[217] = 64'd0;
	mem_0[218] = 64'd0;
	mem_0[219] = 64'd0;
	mem_0[220] = 64'd0;
	mem_0[221] = 64'd0;
	mem_0[222] = 64'd0;
	mem_0[223] = 64'd0;
	mem_0[224] = 64'd0;
	mem_0[225] = 64'd0;
	mem_0[226] = 64'd0;
	mem_0[227] = 64'd0;
	mem_0[228] = 64'd0;
	mem_0[229] = 64'd0;
	mem_0[230] = 64'd0;
	mem_0[231] = 64'd0;
	mem_0[232] = 64'd0;
	mem_0[233] = 64'd0;
	mem_0[234] = 64'd0;
	mem_0[235] = 64'd0;
	mem_0[236] = 64'd0;
	mem_0[237] = 64'd0;
	mem_0[238] = 64'd0;
	mem_0[239] = 64'd0;
	mem_0[240] = 64'd0;
	mem_0[241] = 64'd0;
	mem_0[242] = 64'd0;
	mem_0[243] = 64'd0;
	mem_0[244] = 64'd0;
	mem_0[245] = 64'd0;
	mem_0[246] = 64'd0;
	mem_0[247] = 64'd0;
	mem_0[248] = 64'd0;
	mem_0[249] = 64'd0;
	mem_0[250] = 64'd0;
	mem_0[251] = 64'd0;
	mem_0[252] = 64'd0;
	mem_0[253] = 64'd0;
	mem_0[254] = 64'd0;
	mem_0[255] = 64'd0;
	mem_0[256] = 64'd0;
	mem_0[257] = 64'd0;
	mem_0[258] = 64'd0;
	mem_0[259] = 64'd0;
	mem_0[260] = 64'd0;
	mem_0[261] = 64'd0;
	mem_0[262] = 64'd0;
	mem_0[263] = 64'd0;
	mem_0[264] = 64'd0;
	mem_0[265] = 64'd0;
	mem_0[266] = 64'd0;
	mem_0[267] = 64'd0;
	mem_0[268] = 64'd0;
	mem_0[269] = 64'd0;
	mem_0[270] = 64'd0;
	mem_0[271] = 64'd0;
	mem_0[272] = 64'd0;
	mem_0[273] = 64'd0;
	mem_0[274] = 64'd0;
	mem_0[275] = 64'd0;
	mem_0[276] = 64'd0;
	mem_0[277] = 64'd0;
	mem_0[278] = 64'd0;
	mem_0[279] = 64'd0;
	mem_0[280] = 64'd0;
	mem_0[281] = 64'd0;
	mem_0[282] = 64'd0;
	mem_0[283] = 64'd0;
	mem_0[284] = 64'd0;
	mem_0[285] = 64'd0;
	mem_0[286] = 64'd0;
	mem_0[287] = 64'd0;
	mem_0[288] = 64'd0;
	mem_0[289] = 64'd0;
	mem_0[290] = 64'd0;
	mem_0[291] = 64'd0;
	mem_0[292] = 64'd0;
	mem_0[293] = 64'd0;
	mem_0[294] = 64'd0;
	mem_0[295] = 64'd0;
	mem_0[296] = 64'd0;
	mem_0[297] = 64'd0;
	mem_0[298] = 64'd0;
	mem_0[299] = 64'd0;
	mem_0[300] = 64'd0;
	mem_0[301] = 64'd0;
	mem_0[302] = 64'd0;
	mem_0[303] = 64'd0;
	mem_0[304] = 64'd0;
	mem_0[305] = 64'd0;
	mem_0[306] = 64'd0;
	mem_0[307] = 64'd0;
	mem_0[308] = 64'd0;
	mem_0[309] = 64'd0;
	mem_0[310] = 64'd0;
	mem_0[311] = 64'd0;
	mem_0[312] = 64'd0;
	mem_0[313] = 64'd0;
	mem_0[314] = 64'd0;
	mem_0[315] = 64'd0;
	mem_0[316] = 64'd0;
	mem_0[317] = 64'd0;
	mem_0[318] = 64'd0;
	mem_0[319] = 64'd0;
	mem_0[320] = 64'd0;
	mem_0[321] = 64'd0;
	mem_0[322] = 64'd0;
	mem_0[323] = 64'd0;
	mem_0[324] = 64'd0;
	mem_0[325] = 64'd0;
	mem_0[326] = 64'd0;
	mem_0[327] = 64'd0;
	mem_0[328] = 64'd0;
	mem_0[329] = 64'd0;
	mem_0[330] = 64'd0;
	mem_0[331] = 64'd0;
	mem_0[332] = 64'd0;
	mem_0[333] = 64'd0;
	mem_0[334] = 64'd0;
	mem_0[335] = 64'd0;
	mem_0[336] = 64'd0;
	mem_0[337] = 64'd0;
	mem_0[338] = 64'd0;
	mem_0[339] = 64'd0;
	mem_0[340] = 64'd0;
	mem_0[341] = 64'd0;
	mem_0[342] = 64'd0;
	mem_0[343] = 64'd0;
	mem_0[344] = 64'd0;
	mem_0[345] = 64'd0;
	mem_0[346] = 64'd0;
	mem_0[347] = 64'd0;
	mem_0[348] = 64'd0;
	mem_0[349] = 64'd0;
	mem_0[350] = 64'd0;
	mem_0[351] = 64'd0;
	mem_0[352] = 64'd0;
	mem_0[353] = 64'd0;
	mem_0[354] = 64'd0;
	mem_0[355] = 64'd0;
	mem_0[356] = 64'd0;
	mem_0[357] = 64'd0;
	mem_0[358] = 64'd0;
	mem_0[359] = 64'd0;
	mem_0[360] = 64'd0;
	mem_0[361] = 64'd0;
	mem_0[362] = 64'd0;
	mem_0[363] = 64'd0;
	mem_0[364] = 64'd0;
	mem_0[365] = 64'd0;
	mem_0[366] = 64'd0;
	mem_0[367] = 64'd0;
	mem_0[368] = 64'd0;
	mem_0[369] = 64'd0;
	mem_0[370] = 64'd0;
	mem_0[371] = 64'd0;
	mem_0[372] = 64'd0;
	mem_0[373] = 64'd0;
	mem_0[374] = 64'd0;
	mem_0[375] = 64'd0;
	mem_0[376] = 64'd0;
	mem_0[377] = 64'd0;
	mem_0[378] = 64'd0;
	mem_0[379] = 64'd0;
	mem_0[380] = 64'd0;
	mem_0[381] = 64'd0;
	mem_0[382] = 64'd0;
	mem_0[383] = 64'd0;
	mem_0[384] = 64'd0;
	mem_0[385] = 64'd0;
	mem_0[386] = 64'd0;
	mem_0[387] = 64'd0;
	mem_0[388] = 64'd0;
	mem_0[389] = 64'd0;
	mem_0[390] = 64'd0;
	mem_0[391] = 64'd0;
	mem_0[392] = 64'd0;
	mem_0[393] = 64'd0;
	mem_0[394] = 64'd0;
	mem_0[395] = 64'd0;
	mem_0[396] = 64'd0;
	mem_0[397] = 64'd0;
	mem_0[398] = 64'd0;
	mem_0[399] = 64'd0;
	mem_0[400] = 64'd0;
	mem_0[401] = 64'd0;
	mem_0[402] = 64'd0;
	mem_0[403] = 64'd0;
	mem_0[404] = 64'd0;
	mem_0[405] = 64'd0;
	mem_0[406] = 64'd0;
	mem_0[407] = 64'd0;
	mem_0[408] = 64'd0;
	mem_0[409] = 64'd0;
	mem_0[410] = 64'd0;
	mem_0[411] = 64'd0;
	mem_0[412] = 64'd0;
	mem_0[413] = 64'd0;
	mem_0[414] = 64'd0;
	mem_0[415] = 64'd0;
	mem_0[416] = 64'd0;
	mem_0[417] = 64'd0;
	mem_0[418] = 64'd0;
	mem_0[419] = 64'd0;
	mem_0[420] = 64'd0;
	mem_0[421] = 64'd0;
	mem_0[422] = 64'd0;
	mem_0[423] = 64'd0;
	mem_0[424] = 64'd0;
	mem_0[425] = 64'd0;
	mem_0[426] = 64'd0;
	mem_0[427] = 64'd0;
	mem_0[428] = 64'd0;
	mem_0[429] = 64'd0;
	mem_0[430] = 64'd0;
	mem_0[431] = 64'd0;
	mem_0[432] = 64'd0;
	mem_0[433] = 64'd0;
	mem_0[434] = 64'd0;
	mem_0[435] = 64'd0;
	mem_0[436] = 64'd0;
	mem_0[437] = 64'd0;
	mem_0[438] = 64'd0;
	mem_0[439] = 64'd0;
	mem_0[440] = 64'd0;
	mem_0[441] = 64'd0;
	mem_0[442] = 64'd0;
	mem_0[443] = 64'd0;
	mem_0[444] = 64'd0;
	mem_0[445] = 64'd0;
	mem_0[446] = 64'd0;
	mem_0[447] = 64'd0;
	mem_0[448] = 64'd0;
	mem_0[449] = 64'd0;
	mem_0[450] = 64'd0;
	mem_0[451] = 64'd0;
	mem_0[452] = 64'd0;
	mem_0[453] = 64'd0;
	mem_0[454] = 64'd0;
	mem_0[455] = 64'd0;
	mem_0[456] = 64'd0;
	mem_0[457] = 64'd0;
	mem_0[458] = 64'd0;
	mem_0[459] = 64'd0;
	mem_0[460] = 64'd0;
	mem_0[461] = 64'd0;
	mem_0[462] = 64'd0;
	mem_0[463] = 64'd0;
	mem_0[464] = 64'd0;
	mem_0[465] = 64'd0;
	mem_0[466] = 64'd0;
	mem_0[467] = 64'd0;
	mem_0[468] = 64'd0;
	mem_0[469] = 64'd0;
	mem_0[470] = 64'd0;
	mem_0[471] = 64'd0;
	mem_0[472] = 64'd0;
	mem_0[473] = 64'd0;
	mem_0[474] = 64'd0;
	mem_0[475] = 64'd0;
	mem_0[476] = 64'd0;
	mem_0[477] = 64'd0;
	mem_0[478] = 64'd0;
	mem_0[479] = 64'd0;
	mem_0[480] = 64'd0;
	mem_0[481] = 64'd0;
	mem_0[482] = 64'd0;
	mem_0[483] = 64'd0;
	mem_0[484] = 64'd0;
	mem_0[485] = 64'd0;
	mem_0[486] = 64'd0;
	mem_0[487] = 64'd0;
	mem_0[488] = 64'd0;
	mem_0[489] = 64'd0;
	mem_0[490] = 64'd0;
	mem_0[491] = 64'd0;
	mem_0[492] = 64'd0;
	mem_0[493] = 64'd0;
	mem_0[494] = 64'd0;
	mem_0[495] = 64'd0;
	mem_0[496] = 64'd0;
	mem_0[497] = 64'd0;
	mem_0[498] = 64'd0;
	mem_0[499] = 64'd0;
	mem_0[500] = 64'd0;
	mem_0[501] = 64'd0;
	mem_0[502] = 64'd0;
	mem_0[503] = 64'd0;
	mem_0[504] = 64'd0;
	mem_0[505] = 64'd0;
	mem_0[506] = 64'd0;
	mem_0[507] = 64'd0;
	mem_0[508] = 64'd0;
	mem_0[509] = 64'd0;
	mem_0[510] = 64'd0;
	mem_0[511] = 64'd0;
	mem_0[512] = 64'd0;
	mem_0[513] = 64'd0;
	mem_0[514] = 64'd0;
	mem_0[515] = 64'd0;
	mem_0[516] = 64'd0;
	mem_0[517] = 64'd0;
	mem_0[518] = 64'd0;
	mem_0[519] = 64'd0;
	mem_0[520] = 64'd0;
	mem_0[521] = 64'd0;
	mem_0[522] = 64'd0;
	mem_0[523] = 64'd0;
	mem_0[524] = 64'd0;
	mem_0[525] = 64'd0;
	mem_0[526] = 64'd0;
	mem_0[527] = 64'd0;
	mem_0[528] = 64'd0;
	mem_0[529] = 64'd0;
	mem_0[530] = 64'd0;
	mem_0[531] = 64'd0;
	mem_0[532] = 64'd0;
	mem_0[533] = 64'd0;
	mem_0[534] = 64'd0;
	mem_0[535] = 64'd0;
	mem_0[536] = 64'd0;
	mem_0[537] = 64'd0;
	mem_0[538] = 64'd0;
	mem_0[539] = 64'd0;
	mem_0[540] = 64'd0;
	mem_0[541] = 64'd0;
	mem_0[542] = 64'd0;
	mem_0[543] = 64'd0;
	mem_0[544] = 64'd0;
	mem_0[545] = 64'd0;
	mem_0[546] = 64'd0;
	mem_0[547] = 64'd0;
	mem_0[548] = 64'd0;
	mem_0[549] = 64'd0;
	mem_0[550] = 64'd0;
	mem_0[551] = 64'd0;
	mem_0[552] = 64'd0;
	mem_0[553] = 64'd0;
	mem_0[554] = 64'd0;
	mem_0[555] = 64'd0;
	mem_0[556] = 64'd0;
	mem_0[557] = 64'd0;
	mem_0[558] = 64'd0;
	mem_0[559] = 64'd0;
	mem_0[560] = 64'd0;
	mem_0[561] = 64'd0;
	mem_0[562] = 64'd0;
	mem_0[563] = 64'd0;
	mem_0[564] = 64'd0;
	mem_0[565] = 64'd0;
	mem_0[566] = 64'd0;
	mem_0[567] = 64'd0;
	mem_0[568] = 64'd0;
	mem_0[569] = 64'd0;
	mem_0[570] = 64'd0;
	mem_0[571] = 64'd0;
	mem_0[572] = 64'd0;
	mem_0[573] = 64'd0;
	mem_0[574] = 64'd0;
	mem_0[575] = 64'd0;
	mem_0[576] = 64'd0;
	mem_0[577] = 64'd0;
	mem_0[578] = 64'd0;
	mem_0[579] = 64'd0;
	mem_0[580] = 64'd0;
	mem_0[581] = 64'd0;
	mem_0[582] = 64'd0;
	mem_0[583] = 64'd0;
	mem_0[584] = 64'd0;
	mem_0[585] = 64'd0;
	mem_0[586] = 64'd0;
	mem_0[587] = 64'd0;
	mem_0[588] = 64'd0;
	mem_0[589] = 64'd0;
	mem_0[590] = 64'd0;
	mem_0[591] = 64'd0;
	mem_0[592] = 64'd0;
	mem_0[593] = 64'd0;
	mem_0[594] = 64'd0;
	mem_0[595] = 64'd0;
	mem_0[596] = 64'd0;
	mem_0[597] = 64'd0;
	mem_0[598] = 64'd0;
	mem_0[599] = 64'd0;
	mem_0[600] = 64'd0;
	mem_0[601] = 64'd0;
	mem_0[602] = 64'd0;
	mem_0[603] = 64'd0;
	mem_0[604] = 64'd0;
	mem_0[605] = 64'd0;
	mem_0[606] = 64'd0;
	mem_0[607] = 64'd0;
	mem_0[608] = 64'd0;
	mem_0[609] = 64'd0;
	mem_0[610] = 64'd0;
	mem_0[611] = 64'd0;
	mem_0[612] = 64'd0;
	mem_0[613] = 64'd0;
	mem_0[614] = 64'd0;
	mem_0[615] = 64'd0;
	mem_0[616] = 64'd0;
	mem_0[617] = 64'd0;
	mem_0[618] = 64'd0;
	mem_0[619] = 64'd0;
	mem_0[620] = 64'd0;
	mem_0[621] = 64'd0;
	mem_0[622] = 64'd0;
	mem_0[623] = 64'd0;
	mem_0[624] = 64'd0;
	mem_0[625] = 64'd0;
	mem_0[626] = 64'd0;
	mem_0[627] = 64'd0;
	mem_0[628] = 64'd0;
	mem_0[629] = 64'd0;
	mem_0[630] = 64'd0;
	mem_0[631] = 64'd0;
	mem_0[632] = 64'd0;
	mem_0[633] = 64'd0;
	mem_0[634] = 64'd0;
	mem_0[635] = 64'd0;
	mem_0[636] = 64'd0;
	mem_0[637] = 64'd0;
	mem_0[638] = 64'd0;
	mem_0[639] = 64'd0;
	mem_0[640] = 64'd0;
	mem_0[641] = 64'd0;
	mem_0[642] = 64'd0;
	mem_0[643] = 64'd0;
	mem_0[644] = 64'd0;
	mem_0[645] = 64'd0;
	mem_0[646] = 64'd0;
	mem_0[647] = 64'd0;
	mem_0[648] = 64'd0;
	mem_0[649] = 64'd0;
	mem_0[650] = 64'd0;
	mem_0[651] = 64'd0;
	mem_0[652] = 64'd0;
	mem_0[653] = 64'd0;
	mem_0[654] = 64'd0;
	mem_0[655] = 64'd0;
	mem_0[656] = 64'd0;
	mem_0[657] = 64'd0;
	mem_0[658] = 64'd0;
	mem_0[659] = 64'd0;
	mem_0[660] = 64'd0;
	mem_0[661] = 64'd0;
	mem_0[662] = 64'd0;
	mem_0[663] = 64'd0;
	mem_0[664] = 64'd0;
	mem_0[665] = 64'd0;
	mem_0[666] = 64'd0;
	mem_0[667] = 64'd0;
	mem_0[668] = 64'd0;
	mem_0[669] = 64'd0;
	mem_0[670] = 64'd0;
	mem_0[671] = 64'd0;
	mem_0[672] = 64'd0;
	mem_0[673] = 64'd0;
	mem_0[674] = 64'd0;
	mem_0[675] = 64'd0;
	mem_0[676] = 64'd0;
	mem_0[677] = 64'd0;
	mem_0[678] = 64'd0;
	mem_0[679] = 64'd0;
	mem_0[680] = 64'd0;
	mem_0[681] = 64'd0;
	mem_0[682] = 64'd0;
	mem_0[683] = 64'd0;
	mem_0[684] = 64'd0;
	mem_0[685] = 64'd0;
	mem_0[686] = 64'd0;
	mem_0[687] = 64'd0;
	mem_0[688] = 64'd0;
	mem_0[689] = 64'd0;
	mem_0[690] = 64'd0;
	mem_0[691] = 64'd0;
	mem_0[692] = 64'd0;
	mem_0[693] = 64'd0;
	mem_0[694] = 64'd0;
	mem_0[695] = 64'd0;
	mem_0[696] = 64'd0;
	mem_0[697] = 64'd0;
	mem_0[698] = 64'd0;
	mem_0[699] = 64'd0;
	mem_0[700] = 64'd0;
	mem_0[701] = 64'd0;
	mem_0[702] = 64'd0;
	mem_0[703] = 64'd0;
	mem_0[704] = 64'd0;
	mem_0[705] = 64'd0;
	mem_0[706] = 64'd0;
	mem_0[707] = 64'd0;
	mem_0[708] = 64'd0;
	mem_0[709] = 64'd0;
	mem_0[710] = 64'd0;
	mem_0[711] = 64'd0;
	mem_0[712] = 64'd0;
	mem_0[713] = 64'd0;
	mem_0[714] = 64'd0;
	mem_0[715] = 64'd0;
	mem_0[716] = 64'd0;
	mem_0[717] = 64'd0;
	mem_0[718] = 64'd0;
	mem_0[719] = 64'd0;
	mem_0[720] = 64'd0;
	mem_0[721] = 64'd0;
	mem_0[722] = 64'd0;
	mem_0[723] = 64'd0;
	mem_0[724] = 64'd0;
	mem_0[725] = 64'd0;
	mem_0[726] = 64'd0;
	mem_0[727] = 64'd0;
	mem_0[728] = 64'd0;
	mem_0[729] = 64'd0;
	mem_0[730] = 64'd0;
	mem_0[731] = 64'd0;
	mem_0[732] = 64'd0;
	mem_0[733] = 64'd0;
	mem_0[734] = 64'd0;
	mem_0[735] = 64'd0;
	mem_0[736] = 64'd0;
	mem_0[737] = 64'd0;
	mem_0[738] = 64'd0;
	mem_0[739] = 64'd0;
	mem_0[740] = 64'd0;
	mem_0[741] = 64'd0;
	mem_0[742] = 64'd0;
	mem_0[743] = 64'd0;
	mem_0[744] = 64'd0;
	mem_0[745] = 64'd0;
	mem_0[746] = 64'd0;
	mem_0[747] = 64'd0;
	mem_0[748] = 64'd0;
	mem_0[749] = 64'd0;
	mem_0[750] = 64'd0;
	mem_0[751] = 64'd0;
	mem_0[752] = 64'd0;
	mem_0[753] = 64'd0;
	mem_0[754] = 64'd0;
	mem_0[755] = 64'd0;
	mem_0[756] = 64'd0;
	mem_0[757] = 64'd0;
	mem_0[758] = 64'd0;
	mem_0[759] = 64'd0;
	mem_0[760] = 64'd0;
	mem_0[761] = 64'd0;
	mem_0[762] = 64'd0;
	mem_0[763] = 64'd0;
	mem_0[764] = 64'd0;
	mem_0[765] = 64'd0;
	mem_0[766] = 64'd0;
	mem_0[767] = 64'd0;
	mem_0[768] = 64'd0;
	mem_0[769] = 64'd0;
	mem_0[770] = 64'd0;
	mem_0[771] = 64'd0;
	mem_0[772] = 64'd0;
	mem_0[773] = 64'd0;
	mem_0[774] = 64'd0;
	mem_0[775] = 64'd0;
	mem_0[776] = 64'd0;
	mem_0[777] = 64'd0;
	mem_0[778] = 64'd0;
	mem_0[779] = 64'd0;
	mem_0[780] = 64'd0;
	mem_0[781] = 64'd0;
	mem_0[782] = 64'd0;
	mem_0[783] = 64'd0;
	mem_0[784] = 64'd0;
	mem_0[785] = 64'd0;
	mem_0[786] = 64'd0;
	mem_0[787] = 64'd0;
	mem_0[788] = 64'd0;
	mem_0[789] = 64'd0;
	mem_0[790] = 64'd0;
	mem_0[791] = 64'd0;
	mem_0[792] = 64'd0;
	mem_0[793] = 64'd0;
	mem_0[794] = 64'd0;
	mem_0[795] = 64'd0;
	mem_0[796] = 64'd0;
	mem_0[797] = 64'd0;
	mem_0[798] = 64'd0;
	mem_0[799] = 64'd0;
	mem_0[800] = 64'd0;
	mem_0[801] = 64'd0;
	mem_0[802] = 64'd0;
	mem_0[803] = 64'd0;
	mem_0[804] = 64'd0;
	mem_0[805] = 64'd0;
	mem_0[806] = 64'd0;
	mem_0[807] = 64'd0;
	mem_0[808] = 64'd0;
	mem_0[809] = 64'd0;
	mem_0[810] = 64'd0;
	mem_0[811] = 64'd0;
	mem_0[812] = 64'd0;
	mem_0[813] = 64'd0;
	mem_0[814] = 64'd0;
	mem_0[815] = 64'd0;
	mem_0[816] = 64'd0;
	mem_0[817] = 64'd0;
	mem_0[818] = 64'd0;
	mem_0[819] = 64'd0;
	mem_0[820] = 64'd0;
	mem_0[821] = 64'd0;
	mem_0[822] = 64'd0;
	mem_0[823] = 64'd0;
	mem_0[824] = 64'd0;
	mem_0[825] = 64'd0;
	mem_0[826] = 64'd0;
	mem_0[827] = 64'd0;
	mem_0[828] = 64'd0;
	mem_0[829] = 64'd0;
	mem_0[830] = 64'd0;
	mem_0[831] = 64'd0;
	mem_0[832] = 64'd0;
	mem_0[833] = 64'd0;
	mem_0[834] = 64'd0;
	mem_0[835] = 64'd0;
	mem_0[836] = 64'd0;
	mem_0[837] = 64'd0;
	mem_0[838] = 64'd0;
	mem_0[839] = 64'd0;
	mem_0[840] = 64'd0;
	mem_0[841] = 64'd0;
	mem_0[842] = 64'd0;
	mem_0[843] = 64'd0;
	mem_0[844] = 64'd0;
	mem_0[845] = 64'd0;
	mem_0[846] = 64'd0;
	mem_0[847] = 64'd0;
	mem_0[848] = 64'd0;
	mem_0[849] = 64'd0;
	mem_0[850] = 64'd0;
	mem_0[851] = 64'd0;
	mem_0[852] = 64'd0;
	mem_0[853] = 64'd0;
	mem_0[854] = 64'd0;
	mem_0[855] = 64'd0;
	mem_0[856] = 64'd0;
	mem_0[857] = 64'd0;
	mem_0[858] = 64'd0;
	mem_0[859] = 64'd0;
	mem_0[860] = 64'd0;
	mem_0[861] = 64'd0;
	mem_0[862] = 64'd0;
	mem_0[863] = 64'd0;
	mem_0[864] = 64'd0;
	mem_0[865] = 64'd0;
	mem_0[866] = 64'd0;
	mem_0[867] = 64'd0;
	mem_0[868] = 64'd0;
	mem_0[869] = 64'd0;
	mem_0[870] = 64'd0;
	mem_0[871] = 64'd0;
	mem_0[872] = 64'd0;
	mem_0[873] = 64'd0;
	mem_0[874] = 64'd0;
	mem_0[875] = 64'd0;
	mem_0[876] = 64'd0;
	mem_0[877] = 64'd0;
	mem_0[878] = 64'd0;
	mem_0[879] = 64'd0;
	mem_0[880] = 64'd0;
	mem_0[881] = 64'd0;
	mem_0[882] = 64'd0;
	mem_0[883] = 64'd0;
	mem_0[884] = 64'd0;
	mem_0[885] = 64'd0;
	mem_0[886] = 64'd0;
	mem_0[887] = 64'd0;
	mem_0[888] = 64'd0;
	mem_0[889] = 64'd0;
	mem_0[890] = 64'd0;
	mem_0[891] = 64'd0;
	mem_0[892] = 64'd0;
	mem_0[893] = 64'd0;
	mem_0[894] = 64'd0;
	mem_0[895] = 64'd0;
	mem_0[896] = 64'd0;
	mem_0[897] = 64'd0;
	mem_0[898] = 64'd0;
	mem_0[899] = 64'd0;
	mem_0[900] = 64'd0;
	mem_0[901] = 64'd0;
	mem_0[902] = 64'd0;
	mem_0[903] = 64'd0;
	mem_0[904] = 64'd0;
	mem_0[905] = 64'd0;
	mem_0[906] = 64'd0;
	mem_0[907] = 64'd0;
	mem_0[908] = 64'd0;
	mem_0[909] = 64'd0;
	mem_0[910] = 64'd0;
	mem_0[911] = 64'd0;
	mem_0[912] = 64'd0;
	mem_0[913] = 64'd0;
	mem_0[914] = 64'd0;
	mem_0[915] = 64'd0;
	mem_0[916] = 64'd0;
	mem_0[917] = 64'd0;
	mem_0[918] = 64'd0;
	mem_0[919] = 64'd0;
	mem_0[920] = 64'd0;
	mem_0[921] = 64'd0;
	mem_0[922] = 64'd0;
	mem_0[923] = 64'd0;
	mem_0[924] = 64'd0;
	mem_0[925] = 64'd0;
	mem_0[926] = 64'd0;
	mem_0[927] = 64'd0;
	mem_0[928] = 64'd0;
	mem_0[929] = 64'd0;
	mem_0[930] = 64'd0;
	mem_0[931] = 64'd0;
	mem_0[932] = 64'd0;
	mem_0[933] = 64'd0;
	mem_0[934] = 64'd0;
	mem_0[935] = 64'd0;
	mem_0[936] = 64'd0;
	mem_0[937] = 64'd0;
	mem_0[938] = 64'd0;
	mem_0[939] = 64'd0;
	mem_0[940] = 64'd0;
	mem_0[941] = 64'd0;
	mem_0[942] = 64'd0;
	mem_0[943] = 64'd0;
	mem_0[944] = 64'd0;
	mem_0[945] = 64'd0;
	mem_0[946] = 64'd0;
	mem_0[947] = 64'd0;
	mem_0[948] = 64'd0;
	mem_0[949] = 64'd0;
	mem_0[950] = 64'd0;
	mem_0[951] = 64'd0;
	mem_0[952] = 64'd0;
	mem_0[953] = 64'd0;
	mem_0[954] = 64'd0;
	mem_0[955] = 64'd0;
	mem_0[956] = 64'd0;
	mem_0[957] = 64'd0;
	mem_0[958] = 64'd0;
	mem_0[959] = 64'd0;
	mem_0[960] = 64'd0;
	mem_0[961] = 64'd0;
	mem_0[962] = 64'd0;
	mem_0[963] = 64'd0;
	mem_0[964] = 64'd0;
	mem_0[965] = 64'd0;
	mem_0[966] = 64'd0;
	mem_0[967] = 64'd0;
	mem_0[968] = 64'd0;
	mem_0[969] = 64'd0;
	mem_0[970] = 64'd0;
	mem_0[971] = 64'd0;
	mem_0[972] = 64'd0;
	mem_0[973] = 64'd0;
	mem_0[974] = 64'd0;
	mem_0[975] = 64'd0;
	mem_0[976] = 64'd0;
	mem_0[977] = 64'd0;
	mem_0[978] = 64'd0;
	mem_0[979] = 64'd0;
	mem_0[980] = 64'd0;
	mem_0[981] = 64'd0;
	mem_0[982] = 64'd0;
	mem_0[983] = 64'd0;
	mem_0[984] = 64'd0;
	mem_0[985] = 64'd0;
	mem_0[986] = 64'd0;
	mem_0[987] = 64'd0;
	mem_0[988] = 64'd0;
	mem_0[989] = 64'd0;
	mem_0[990] = 64'd0;
	mem_0[991] = 64'd0;
	mem_0[992] = 64'd0;
	mem_0[993] = 64'd0;
	mem_0[994] = 64'd0;
	mem_0[995] = 64'd0;
	mem_0[996] = 64'd0;
	mem_0[997] = 64'd0;
	mem_0[998] = 64'd0;
	mem_0[999] = 64'd0;
	mem_0[1000] = 64'd0;
	mem_0[1001] = 64'd0;
	mem_0[1002] = 64'd0;
	mem_0[1003] = 64'd0;
	mem_0[1004] = 64'd0;
	mem_0[1005] = 64'd0;
	mem_0[1006] = 64'd0;
	mem_0[1007] = 64'd0;
	mem_0[1008] = 64'd0;
	mem_0[1009] = 64'd0;
	mem_0[1010] = 64'd0;
	mem_0[1011] = 64'd0;
	mem_0[1012] = 64'd0;
	mem_0[1013] = 64'd0;
	mem_0[1014] = 64'd0;
	mem_0[1015] = 64'd0;
	mem_0[1016] = 64'd0;
	mem_0[1017] = 64'd0;
	mem_0[1018] = 64'd0;
	mem_0[1019] = 64'd0;
	mem_0[1020] = 64'd0;
	mem_0[1021] = 64'd0;
	mem_0[1022] = 64'd0;
	mem_0[1023] = 64'd0;
	mem_1[0] = 64'd0;
	mem_1[1] = 64'd0;
	mem_1[2] = 64'd0;
	mem_1[3] = 64'd0;
	mem_1[4] = 64'd0;
	mem_1[5] = 64'd0;
	mem_1[6] = 64'd0;
	mem_1[7] = 64'd0;
	mem_1[8] = 64'd0;
	mem_1[9] = 64'd0;
	mem_1[10] = 64'd0;
	mem_1[11] = 64'd0;
	mem_1[12] = 64'd0;
	mem_1[13] = 64'd0;
	mem_1[14] = 64'd0;
	mem_1[15] = 64'd0;
	mem_1[16] = 64'd0;
	mem_1[17] = 64'd0;
	mem_1[18] = 64'd0;
	mem_1[19] = 64'd0;
	mem_1[20] = 64'd0;
	mem_1[21] = 64'd0;
	mem_1[22] = 64'd0;
	mem_1[23] = 64'd0;
	mem_1[24] = 64'd0;
	mem_1[25] = 64'd0;
	mem_1[26] = 64'd0;
	mem_1[27] = 64'd0;
	mem_1[28] = 64'd0;
	mem_1[29] = 64'd0;
	mem_1[30] = 64'd0;
	mem_1[31] = 64'd0;
	mem_1[32] = 64'd0;
	mem_1[33] = 64'd0;
	mem_1[34] = 64'd0;
	mem_1[35] = 64'd0;
	mem_1[36] = 64'd0;
	mem_1[37] = 64'd0;
	mem_1[38] = 64'd0;
	mem_1[39] = 64'd0;
	mem_1[40] = 64'd0;
	mem_1[41] = 64'd0;
	mem_1[42] = 64'd0;
	mem_1[43] = 64'd0;
	mem_1[44] = 64'd0;
	mem_1[45] = 64'd0;
	mem_1[46] = 64'd0;
	mem_1[47] = 64'd0;
	mem_1[48] = 64'd0;
	mem_1[49] = 64'd0;
	mem_1[50] = 64'd0;
	mem_1[51] = 64'd0;
	mem_1[52] = 64'd0;
	mem_1[53] = 64'd0;
	mem_1[54] = 64'd0;
	mem_1[55] = 64'd0;
	mem_1[56] = 64'd0;
	mem_1[57] = 64'd0;
	mem_1[58] = 64'd0;
	mem_1[59] = 64'd0;
	mem_1[60] = 64'd0;
	mem_1[61] = 64'd0;
	mem_1[62] = 64'd0;
	mem_1[63] = 64'd0;
	mem_1[64] = 64'd0;
	mem_1[65] = 64'd0;
	mem_1[66] = 64'd0;
	mem_1[67] = 64'd0;
	mem_1[68] = 64'd0;
	mem_1[69] = 64'd0;
	mem_1[70] = 64'd0;
	mem_1[71] = 64'd0;
	mem_1[72] = 64'd0;
	mem_1[73] = 64'd0;
	mem_1[74] = 64'd0;
	mem_1[75] = 64'd0;
	mem_1[76] = 64'd0;
	mem_1[77] = 64'd0;
	mem_1[78] = 64'd0;
	mem_1[79] = 64'd0;
	mem_1[80] = 64'd0;
	mem_1[81] = 64'd0;
	mem_1[82] = 64'd0;
	mem_1[83] = 64'd0;
	mem_1[84] = 64'd0;
	mem_1[85] = 64'd0;
	mem_1[86] = 64'd0;
	mem_1[87] = 64'd0;
	mem_1[88] = 64'd0;
	mem_1[89] = 64'd0;
	mem_1[90] = 64'd0;
	mem_1[91] = 64'd0;
	mem_1[92] = 64'd0;
	mem_1[93] = 64'd0;
	mem_1[94] = 64'd0;
	mem_1[95] = 64'd0;
	mem_1[96] = 64'd0;
	mem_1[97] = 64'd0;
	mem_1[98] = 64'd0;
	mem_1[99] = 64'd0;
	mem_1[100] = 64'd0;
	mem_1[101] = 64'd0;
	mem_1[102] = 64'd0;
	mem_1[103] = 64'd0;
	mem_1[104] = 64'd0;
	mem_1[105] = 64'd0;
	mem_1[106] = 64'd0;
	mem_1[107] = 64'd0;
	mem_1[108] = 64'd0;
	mem_1[109] = 64'd0;
	mem_1[110] = 64'd0;
	mem_1[111] = 64'd0;
	mem_1[112] = 64'd0;
	mem_1[113] = 64'd0;
	mem_1[114] = 64'd0;
	mem_1[115] = 64'd0;
	mem_1[116] = 64'd0;
	mem_1[117] = 64'd0;
	mem_1[118] = 64'd0;
	mem_1[119] = 64'd0;
	mem_1[120] = 64'd0;
	mem_1[121] = 64'd0;
	mem_1[122] = 64'd0;
	mem_1[123] = 64'd0;
	mem_1[124] = 64'd0;
	mem_1[125] = 64'd0;
	mem_1[126] = 64'd0;
	mem_1[127] = 64'd0;
	mem_1[128] = 64'd0;
	mem_1[129] = 64'd0;
	mem_1[130] = 64'd0;
	mem_1[131] = 64'd0;
	mem_1[132] = 64'd0;
	mem_1[133] = 64'd0;
	mem_1[134] = 64'd0;
	mem_1[135] = 64'd0;
	mem_1[136] = 64'd0;
	mem_1[137] = 64'd0;
	mem_1[138] = 64'd0;
	mem_1[139] = 64'd0;
	mem_1[140] = 64'd0;
	mem_1[141] = 64'd0;
	mem_1[142] = 64'd0;
	mem_1[143] = 64'd0;
	mem_1[144] = 64'd0;
	mem_1[145] = 64'd0;
	mem_1[146] = 64'd0;
	mem_1[147] = 64'd0;
	mem_1[148] = 64'd0;
	mem_1[149] = 64'd0;
	mem_1[150] = 64'd0;
	mem_1[151] = 64'd0;
	mem_1[152] = 64'd0;
	mem_1[153] = 64'd0;
	mem_1[154] = 64'd0;
	mem_1[155] = 64'd0;
	mem_1[156] = 64'd0;
	mem_1[157] = 64'd0;
	mem_1[158] = 64'd0;
	mem_1[159] = 64'd0;
	mem_1[160] = 64'd0;
	mem_1[161] = 64'd0;
	mem_1[162] = 64'd0;
	mem_1[163] = 64'd0;
	mem_1[164] = 64'd0;
	mem_1[165] = 64'd0;
	mem_1[166] = 64'd0;
	mem_1[167] = 64'd0;
	mem_1[168] = 64'd0;
	mem_1[169] = 64'd0;
	mem_1[170] = 64'd0;
	mem_1[171] = 64'd0;
	mem_1[172] = 64'd0;
	mem_1[173] = 64'd0;
	mem_1[174] = 64'd0;
	mem_1[175] = 64'd0;
	mem_1[176] = 64'd0;
	mem_1[177] = 64'd0;
	mem_1[178] = 64'd0;
	mem_1[179] = 64'd0;
	mem_1[180] = 64'd0;
	mem_1[181] = 64'd0;
	mem_1[182] = 64'd0;
	mem_1[183] = 64'd0;
	mem_1[184] = 64'd0;
	mem_1[185] = 64'd0;
	mem_1[186] = 64'd0;
	mem_1[187] = 64'd0;
	mem_1[188] = 64'd0;
	mem_1[189] = 64'd0;
	mem_1[190] = 64'd0;
	mem_1[191] = 64'd0;
	mem_1[192] = 64'd0;
	mem_1[193] = 64'd0;
	mem_1[194] = 64'd0;
	mem_1[195] = 64'd0;
	mem_1[196] = 64'd0;
	mem_1[197] = 64'd0;
	mem_1[198] = 64'd0;
	mem_1[199] = 64'd0;
	mem_1[200] = 64'd0;
	mem_1[201] = 64'd0;
	mem_1[202] = 64'd0;
	mem_1[203] = 64'd0;
	mem_1[204] = 64'd0;
	mem_1[205] = 64'd0;
	mem_1[206] = 64'd0;
	mem_1[207] = 64'd0;
	mem_1[208] = 64'd0;
	mem_1[209] = 64'd0;
	mem_1[210] = 64'd0;
	mem_1[211] = 64'd0;
	mem_1[212] = 64'd0;
	mem_1[213] = 64'd0;
	mem_1[214] = 64'd0;
	mem_1[215] = 64'd0;
	mem_1[216] = 64'd0;
	mem_1[217] = 64'd0;
	mem_1[218] = 64'd0;
	mem_1[219] = 64'd0;
	mem_1[220] = 64'd0;
	mem_1[221] = 64'd0;
	mem_1[222] = 64'd0;
	mem_1[223] = 64'd0;
	mem_1[224] = 64'd0;
	mem_1[225] = 64'd0;
	mem_1[226] = 64'd0;
	mem_1[227] = 64'd0;
	mem_1[228] = 64'd0;
	mem_1[229] = 64'd0;
	mem_1[230] = 64'd0;
	mem_1[231] = 64'd0;
	mem_1[232] = 64'd0;
	mem_1[233] = 64'd0;
	mem_1[234] = 64'd0;
	mem_1[235] = 64'd0;
	mem_1[236] = 64'd0;
	mem_1[237] = 64'd0;
	mem_1[238] = 64'd0;
	mem_1[239] = 64'd0;
	mem_1[240] = 64'd0;
	mem_1[241] = 64'd0;
	mem_1[242] = 64'd0;
	mem_1[243] = 64'd0;
	mem_1[244] = 64'd0;
	mem_1[245] = 64'd0;
	mem_1[246] = 64'd0;
	mem_1[247] = 64'd0;
	mem_1[248] = 64'd0;
	mem_1[249] = 64'd0;
	mem_1[250] = 64'd0;
	mem_1[251] = 64'd0;
	mem_1[252] = 64'd0;
	mem_1[253] = 64'd0;
	mem_1[254] = 64'd0;
	mem_1[255] = 64'd0;
	mem_1[256] = 64'd0;
	mem_1[257] = 64'd0;
	mem_1[258] = 64'd0;
	mem_1[259] = 64'd0;
	mem_1[260] = 64'd0;
	mem_1[261] = 64'd0;
	mem_1[262] = 64'd0;
	mem_1[263] = 64'd0;
	mem_1[264] = 64'd0;
	mem_1[265] = 64'd0;
	mem_1[266] = 64'd0;
	mem_1[267] = 64'd0;
	mem_1[268] = 64'd0;
	mem_1[269] = 64'd0;
	mem_1[270] = 64'd0;
	mem_1[271] = 64'd0;
	mem_1[272] = 64'd0;
	mem_1[273] = 64'd0;
	mem_1[274] = 64'd0;
	mem_1[275] = 64'd0;
	mem_1[276] = 64'd0;
	mem_1[277] = 64'd0;
	mem_1[278] = 64'd0;
	mem_1[279] = 64'd0;
	mem_1[280] = 64'd0;
	mem_1[281] = 64'd0;
	mem_1[282] = 64'd0;
	mem_1[283] = 64'd0;
	mem_1[284] = 64'd0;
	mem_1[285] = 64'd0;
	mem_1[286] = 64'd0;
	mem_1[287] = 64'd0;
	mem_1[288] = 64'd0;
	mem_1[289] = 64'd0;
	mem_1[290] = 64'd0;
	mem_1[291] = 64'd0;
	mem_1[292] = 64'd0;
	mem_1[293] = 64'd0;
	mem_1[294] = 64'd0;
	mem_1[295] = 64'd0;
	mem_1[296] = 64'd0;
	mem_1[297] = 64'd0;
	mem_1[298] = 64'd0;
	mem_1[299] = 64'd0;
	mem_1[300] = 64'd0;
	mem_1[301] = 64'd0;
	mem_1[302] = 64'd0;
	mem_1[303] = 64'd0;
	mem_1[304] = 64'd0;
	mem_1[305] = 64'd0;
	mem_1[306] = 64'd0;
	mem_1[307] = 64'd0;
	mem_1[308] = 64'd0;
	mem_1[309] = 64'd0;
	mem_1[310] = 64'd0;
	mem_1[311] = 64'd0;
	mem_1[312] = 64'd0;
	mem_1[313] = 64'd0;
	mem_1[314] = 64'd0;
	mem_1[315] = 64'd0;
	mem_1[316] = 64'd0;
	mem_1[317] = 64'd0;
	mem_1[318] = 64'd0;
	mem_1[319] = 64'd0;
	mem_1[320] = 64'd0;
	mem_1[321] = 64'd0;
	mem_1[322] = 64'd0;
	mem_1[323] = 64'd0;
	mem_1[324] = 64'd0;
	mem_1[325] = 64'd0;
	mem_1[326] = 64'd0;
	mem_1[327] = 64'd0;
	mem_1[328] = 64'd0;
	mem_1[329] = 64'd0;
	mem_1[330] = 64'd0;
	mem_1[331] = 64'd0;
	mem_1[332] = 64'd0;
	mem_1[333] = 64'd0;
	mem_1[334] = 64'd0;
	mem_1[335] = 64'd0;
	mem_1[336] = 64'd0;
	mem_1[337] = 64'd0;
	mem_1[338] = 64'd0;
	mem_1[339] = 64'd0;
	mem_1[340] = 64'd0;
	mem_1[341] = 64'd0;
	mem_1[342] = 64'd0;
	mem_1[343] = 64'd0;
	mem_1[344] = 64'd0;
	mem_1[345] = 64'd0;
	mem_1[346] = 64'd0;
	mem_1[347] = 64'd0;
	mem_1[348] = 64'd0;
	mem_1[349] = 64'd0;
	mem_1[350] = 64'd0;
	mem_1[351] = 64'd0;
	mem_1[352] = 64'd0;
	mem_1[353] = 64'd0;
	mem_1[354] = 64'd0;
	mem_1[355] = 64'd0;
	mem_1[356] = 64'd0;
	mem_1[357] = 64'd0;
	mem_1[358] = 64'd0;
	mem_1[359] = 64'd0;
	mem_1[360] = 64'd0;
	mem_1[361] = 64'd0;
	mem_1[362] = 64'd0;
	mem_1[363] = 64'd0;
	mem_1[364] = 64'd0;
	mem_1[365] = 64'd0;
	mem_1[366] = 64'd0;
	mem_1[367] = 64'd0;
	mem_1[368] = 64'd0;
	mem_1[369] = 64'd0;
	mem_1[370] = 64'd0;
	mem_1[371] = 64'd0;
	mem_1[372] = 64'd0;
	mem_1[373] = 64'd0;
	mem_1[374] = 64'd0;
	mem_1[375] = 64'd0;
	mem_1[376] = 64'd0;
	mem_1[377] = 64'd0;
	mem_1[378] = 64'd0;
	mem_1[379] = 64'd0;
	mem_1[380] = 64'd0;
	mem_1[381] = 64'd0;
	mem_1[382] = 64'd0;
	mem_1[383] = 64'd0;
	mem_1[384] = 64'd0;
	mem_1[385] = 64'd0;
	mem_1[386] = 64'd0;
	mem_1[387] = 64'd0;
	mem_1[388] = 64'd0;
	mem_1[389] = 64'd0;
	mem_1[390] = 64'd0;
	mem_1[391] = 64'd0;
	mem_1[392] = 64'd0;
	mem_1[393] = 64'd0;
	mem_1[394] = 64'd0;
	mem_1[395] = 64'd0;
	mem_1[396] = 64'd0;
	mem_1[397] = 64'd0;
	mem_1[398] = 64'd0;
	mem_1[399] = 64'd0;
	mem_1[400] = 64'd0;
	mem_1[401] = 64'd0;
	mem_1[402] = 64'd0;
	mem_1[403] = 64'd0;
	mem_1[404] = 64'd0;
	mem_1[405] = 64'd0;
	mem_1[406] = 64'd0;
	mem_1[407] = 64'd0;
	mem_1[408] = 64'd0;
	mem_1[409] = 64'd0;
	mem_1[410] = 64'd0;
	mem_1[411] = 64'd0;
	mem_1[412] = 64'd0;
	mem_1[413] = 64'd0;
	mem_1[414] = 64'd0;
	mem_1[415] = 64'd0;
	mem_1[416] = 64'd0;
	mem_1[417] = 64'd0;
	mem_1[418] = 64'd0;
	mem_1[419] = 64'd0;
	mem_1[420] = 64'd0;
	mem_1[421] = 64'd0;
	mem_1[422] = 64'd0;
	mem_1[423] = 64'd0;
	mem_1[424] = 64'd0;
	mem_1[425] = 64'd0;
	mem_1[426] = 64'd0;
	mem_1[427] = 64'd0;
	mem_1[428] = 64'd0;
	mem_1[429] = 64'd0;
	mem_1[430] = 64'd0;
	mem_1[431] = 64'd0;
	mem_1[432] = 64'd0;
	mem_1[433] = 64'd0;
	mem_1[434] = 64'd0;
	mem_1[435] = 64'd0;
	mem_1[436] = 64'd0;
	mem_1[437] = 64'd0;
	mem_1[438] = 64'd0;
	mem_1[439] = 64'd0;
	mem_1[440] = 64'd0;
	mem_1[441] = 64'd0;
	mem_1[442] = 64'd0;
	mem_1[443] = 64'd0;
	mem_1[444] = 64'd0;
	mem_1[445] = 64'd0;
	mem_1[446] = 64'd0;
	mem_1[447] = 64'd0;
	mem_1[448] = 64'd0;
	mem_1[449] = 64'd0;
	mem_1[450] = 64'd0;
	mem_1[451] = 64'd0;
	mem_1[452] = 64'd0;
	mem_1[453] = 64'd0;
	mem_1[454] = 64'd0;
	mem_1[455] = 64'd0;
	mem_1[456] = 64'd0;
	mem_1[457] = 64'd0;
	mem_1[458] = 64'd0;
	mem_1[459] = 64'd0;
	mem_1[460] = 64'd0;
	mem_1[461] = 64'd0;
	mem_1[462] = 64'd0;
	mem_1[463] = 64'd0;
	mem_1[464] = 64'd0;
	mem_1[465] = 64'd0;
	mem_1[466] = 64'd0;
	mem_1[467] = 64'd0;
	mem_1[468] = 64'd0;
	mem_1[469] = 64'd0;
	mem_1[470] = 64'd0;
	mem_1[471] = 64'd0;
	mem_1[472] = 64'd0;
	mem_1[473] = 64'd0;
	mem_1[474] = 64'd0;
	mem_1[475] = 64'd0;
	mem_1[476] = 64'd0;
	mem_1[477] = 64'd0;
	mem_1[478] = 64'd0;
	mem_1[479] = 64'd0;
	mem_1[480] = 64'd0;
	mem_1[481] = 64'd0;
	mem_1[482] = 64'd0;
	mem_1[483] = 64'd0;
	mem_1[484] = 64'd0;
	mem_1[485] = 64'd0;
	mem_1[486] = 64'd0;
	mem_1[487] = 64'd0;
	mem_1[488] = 64'd0;
	mem_1[489] = 64'd0;
	mem_1[490] = 64'd0;
	mem_1[491] = 64'd0;
	mem_1[492] = 64'd0;
	mem_1[493] = 64'd0;
	mem_1[494] = 64'd0;
	mem_1[495] = 64'd0;
	mem_1[496] = 64'd0;
	mem_1[497] = 64'd0;
	mem_1[498] = 64'd0;
	mem_1[499] = 64'd0;
	mem_1[500] = 64'd0;
	mem_1[501] = 64'd0;
	mem_1[502] = 64'd0;
	mem_1[503] = 64'd0;
	mem_1[504] = 64'd0;
	mem_1[505] = 64'd0;
	mem_1[506] = 64'd0;
	mem_1[507] = 64'd0;
	mem_1[508] = 64'd0;
	mem_1[509] = 64'd0;
	mem_1[510] = 64'd0;
	mem_1[511] = 64'd0;
	mem_1[512] = 64'd0;
	mem_1[513] = 64'd0;
	mem_1[514] = 64'd0;
	mem_1[515] = 64'd0;
	mem_1[516] = 64'd0;
	mem_1[517] = 64'd0;
	mem_1[518] = 64'd0;
	mem_1[519] = 64'd0;
	mem_1[520] = 64'd0;
	mem_1[521] = 64'd0;
	mem_1[522] = 64'd0;
	mem_1[523] = 64'd0;
	mem_1[524] = 64'd0;
	mem_1[525] = 64'd0;
	mem_1[526] = 64'd0;
	mem_1[527] = 64'd0;
	mem_1[528] = 64'd0;
	mem_1[529] = 64'd0;
	mem_1[530] = 64'd0;
	mem_1[531] = 64'd0;
	mem_1[532] = 64'd0;
	mem_1[533] = 64'd0;
	mem_1[534] = 64'd0;
	mem_1[535] = 64'd0;
	mem_1[536] = 64'd0;
	mem_1[537] = 64'd0;
	mem_1[538] = 64'd0;
	mem_1[539] = 64'd0;
	mem_1[540] = 64'd0;
	mem_1[541] = 64'd0;
	mem_1[542] = 64'd0;
	mem_1[543] = 64'd0;
	mem_1[544] = 64'd0;
	mem_1[545] = 64'd0;
	mem_1[546] = 64'd0;
	mem_1[547] = 64'd0;
	mem_1[548] = 64'd0;
	mem_1[549] = 64'd0;
	mem_1[550] = 64'd0;
	mem_1[551] = 64'd0;
	mem_1[552] = 64'd0;
	mem_1[553] = 64'd0;
	mem_1[554] = 64'd0;
	mem_1[555] = 64'd0;
	mem_1[556] = 64'd0;
	mem_1[557] = 64'd0;
	mem_1[558] = 64'd0;
	mem_1[559] = 64'd0;
	mem_1[560] = 64'd0;
	mem_1[561] = 64'd0;
	mem_1[562] = 64'd0;
	mem_1[563] = 64'd0;
	mem_1[564] = 64'd0;
	mem_1[565] = 64'd0;
	mem_1[566] = 64'd0;
	mem_1[567] = 64'd0;
	mem_1[568] = 64'd0;
	mem_1[569] = 64'd0;
	mem_1[570] = 64'd0;
	mem_1[571] = 64'd0;
	mem_1[572] = 64'd0;
	mem_1[573] = 64'd0;
	mem_1[574] = 64'd0;
	mem_1[575] = 64'd0;
	mem_1[576] = 64'd0;
	mem_1[577] = 64'd0;
	mem_1[578] = 64'd0;
	mem_1[579] = 64'd0;
	mem_1[580] = 64'd0;
	mem_1[581] = 64'd0;
	mem_1[582] = 64'd0;
	mem_1[583] = 64'd0;
	mem_1[584] = 64'd0;
	mem_1[585] = 64'd0;
	mem_1[586] = 64'd0;
	mem_1[587] = 64'd0;
	mem_1[588] = 64'd0;
	mem_1[589] = 64'd0;
	mem_1[590] = 64'd0;
	mem_1[591] = 64'd0;
	mem_1[592] = 64'd0;
	mem_1[593] = 64'd0;
	mem_1[594] = 64'd0;
	mem_1[595] = 64'd0;
	mem_1[596] = 64'd0;
	mem_1[597] = 64'd0;
	mem_1[598] = 64'd0;
	mem_1[599] = 64'd0;
	mem_1[600] = 64'd0;
	mem_1[601] = 64'd0;
	mem_1[602] = 64'd0;
	mem_1[603] = 64'd0;
	mem_1[604] = 64'd0;
	mem_1[605] = 64'd0;
	mem_1[606] = 64'd0;
	mem_1[607] = 64'd0;
	mem_1[608] = 64'd0;
	mem_1[609] = 64'd0;
	mem_1[610] = 64'd0;
	mem_1[611] = 64'd0;
	mem_1[612] = 64'd0;
	mem_1[613] = 64'd0;
	mem_1[614] = 64'd0;
	mem_1[615] = 64'd0;
	mem_1[616] = 64'd0;
	mem_1[617] = 64'd0;
	mem_1[618] = 64'd0;
	mem_1[619] = 64'd0;
	mem_1[620] = 64'd0;
	mem_1[621] = 64'd0;
	mem_1[622] = 64'd0;
	mem_1[623] = 64'd0;
	mem_1[624] = 64'd0;
	mem_1[625] = 64'd0;
	mem_1[626] = 64'd0;
	mem_1[627] = 64'd0;
	mem_1[628] = 64'd0;
	mem_1[629] = 64'd0;
	mem_1[630] = 64'd0;
	mem_1[631] = 64'd0;
	mem_1[632] = 64'd0;
	mem_1[633] = 64'd0;
	mem_1[634] = 64'd0;
	mem_1[635] = 64'd0;
	mem_1[636] = 64'd0;
	mem_1[637] = 64'd0;
	mem_1[638] = 64'd0;
	mem_1[639] = 64'd0;
	mem_1[640] = 64'd0;
	mem_1[641] = 64'd0;
	mem_1[642] = 64'd0;
	mem_1[643] = 64'd0;
	mem_1[644] = 64'd0;
	mem_1[645] = 64'd0;
	mem_1[646] = 64'd0;
	mem_1[647] = 64'd0;
	mem_1[648] = 64'd0;
	mem_1[649] = 64'd0;
	mem_1[650] = 64'd0;
	mem_1[651] = 64'd0;
	mem_1[652] = 64'd0;
	mem_1[653] = 64'd0;
	mem_1[654] = 64'd0;
	mem_1[655] = 64'd0;
	mem_1[656] = 64'd0;
	mem_1[657] = 64'd0;
	mem_1[658] = 64'd0;
	mem_1[659] = 64'd0;
	mem_1[660] = 64'd0;
	mem_1[661] = 64'd0;
	mem_1[662] = 64'd0;
	mem_1[663] = 64'd0;
	mem_1[664] = 64'd0;
	mem_1[665] = 64'd0;
	mem_1[666] = 64'd0;
	mem_1[667] = 64'd0;
	mem_1[668] = 64'd0;
	mem_1[669] = 64'd0;
	mem_1[670] = 64'd0;
	mem_1[671] = 64'd0;
	mem_1[672] = 64'd0;
	mem_1[673] = 64'd0;
	mem_1[674] = 64'd0;
	mem_1[675] = 64'd0;
	mem_1[676] = 64'd0;
	mem_1[677] = 64'd0;
	mem_1[678] = 64'd0;
	mem_1[679] = 64'd0;
	mem_1[680] = 64'd0;
	mem_1[681] = 64'd0;
	mem_1[682] = 64'd0;
	mem_1[683] = 64'd0;
	mem_1[684] = 64'd0;
	mem_1[685] = 64'd0;
	mem_1[686] = 64'd0;
	mem_1[687] = 64'd0;
	mem_1[688] = 64'd0;
	mem_1[689] = 64'd0;
	mem_1[690] = 64'd0;
	mem_1[691] = 64'd0;
	mem_1[692] = 64'd0;
	mem_1[693] = 64'd0;
	mem_1[694] = 64'd0;
	mem_1[695] = 64'd0;
	mem_1[696] = 64'd0;
	mem_1[697] = 64'd0;
	mem_1[698] = 64'd0;
	mem_1[699] = 64'd0;
	mem_1[700] = 64'd0;
	mem_1[701] = 64'd0;
	mem_1[702] = 64'd0;
	mem_1[703] = 64'd0;
	mem_1[704] = 64'd0;
	mem_1[705] = 64'd0;
	mem_1[706] = 64'd0;
	mem_1[707] = 64'd0;
	mem_1[708] = 64'd0;
	mem_1[709] = 64'd0;
	mem_1[710] = 64'd0;
	mem_1[711] = 64'd0;
	mem_1[712] = 64'd0;
	mem_1[713] = 64'd0;
	mem_1[714] = 64'd0;
	mem_1[715] = 64'd0;
	mem_1[716] = 64'd0;
	mem_1[717] = 64'd0;
	mem_1[718] = 64'd0;
	mem_1[719] = 64'd0;
	mem_1[720] = 64'd0;
	mem_1[721] = 64'd0;
	mem_1[722] = 64'd0;
	mem_1[723] = 64'd0;
	mem_1[724] = 64'd0;
	mem_1[725] = 64'd0;
	mem_1[726] = 64'd0;
	mem_1[727] = 64'd0;
	mem_1[728] = 64'd0;
	mem_1[729] = 64'd0;
	mem_1[730] = 64'd0;
	mem_1[731] = 64'd0;
	mem_1[732] = 64'd0;
	mem_1[733] = 64'd0;
	mem_1[734] = 64'd0;
	mem_1[735] = 64'd0;
	mem_1[736] = 64'd0;
	mem_1[737] = 64'd0;
	mem_1[738] = 64'd0;
	mem_1[739] = 64'd0;
	mem_1[740] = 64'd0;
	mem_1[741] = 64'd0;
	mem_1[742] = 64'd0;
	mem_1[743] = 64'd0;
	mem_1[744] = 64'd0;
	mem_1[745] = 64'd0;
	mem_1[746] = 64'd0;
	mem_1[747] = 64'd0;
	mem_1[748] = 64'd0;
	mem_1[749] = 64'd0;
	mem_1[750] = 64'd0;
	mem_1[751] = 64'd0;
	mem_1[752] = 64'd0;
	mem_1[753] = 64'd0;
	mem_1[754] = 64'd0;
	mem_1[755] = 64'd0;
	mem_1[756] = 64'd0;
	mem_1[757] = 64'd0;
	mem_1[758] = 64'd0;
	mem_1[759] = 64'd0;
	mem_1[760] = 64'd0;
	mem_1[761] = 64'd0;
	mem_1[762] = 64'd0;
	mem_1[763] = 64'd0;
	mem_1[764] = 64'd0;
	mem_1[765] = 64'd0;
	mem_1[766] = 64'd0;
	mem_1[767] = 64'd0;
	mem_1[768] = 64'd0;
	mem_1[769] = 64'd0;
	mem_1[770] = 64'd0;
	mem_1[771] = 64'd0;
	mem_1[772] = 64'd0;
	mem_1[773] = 64'd0;
	mem_1[774] = 64'd0;
	mem_1[775] = 64'd0;
	mem_1[776] = 64'd0;
	mem_1[777] = 64'd0;
	mem_1[778] = 64'd0;
	mem_1[779] = 64'd0;
	mem_1[780] = 64'd0;
	mem_1[781] = 64'd0;
	mem_1[782] = 64'd0;
	mem_1[783] = 64'd0;
	mem_1[784] = 64'd0;
	mem_1[785] = 64'd0;
	mem_1[786] = 64'd0;
	mem_1[787] = 64'd0;
	mem_1[788] = 64'd0;
	mem_1[789] = 64'd0;
	mem_1[790] = 64'd0;
	mem_1[791] = 64'd0;
	mem_1[792] = 64'd0;
	mem_1[793] = 64'd0;
	mem_1[794] = 64'd0;
	mem_1[795] = 64'd0;
	mem_1[796] = 64'd0;
	mem_1[797] = 64'd0;
	mem_1[798] = 64'd0;
	mem_1[799] = 64'd0;
	mem_1[800] = 64'd0;
	mem_1[801] = 64'd0;
	mem_1[802] = 64'd0;
	mem_1[803] = 64'd0;
	mem_1[804] = 64'd0;
	mem_1[805] = 64'd0;
	mem_1[806] = 64'd0;
	mem_1[807] = 64'd0;
	mem_1[808] = 64'd0;
	mem_1[809] = 64'd0;
	mem_1[810] = 64'd0;
	mem_1[811] = 64'd0;
	mem_1[812] = 64'd0;
	mem_1[813] = 64'd0;
	mem_1[814] = 64'd0;
	mem_1[815] = 64'd0;
	mem_1[816] = 64'd0;
	mem_1[817] = 64'd0;
	mem_1[818] = 64'd0;
	mem_1[819] = 64'd0;
	mem_1[820] = 64'd0;
	mem_1[821] = 64'd0;
	mem_1[822] = 64'd0;
	mem_1[823] = 64'd0;
	mem_1[824] = 64'd0;
	mem_1[825] = 64'd0;
	mem_1[826] = 64'd0;
	mem_1[827] = 64'd0;
	mem_1[828] = 64'd0;
	mem_1[829] = 64'd0;
	mem_1[830] = 64'd0;
	mem_1[831] = 64'd0;
	mem_1[832] = 64'd0;
	mem_1[833] = 64'd0;
	mem_1[834] = 64'd0;
	mem_1[835] = 64'd0;
	mem_1[836] = 64'd0;
	mem_1[837] = 64'd0;
	mem_1[838] = 64'd0;
	mem_1[839] = 64'd0;
	mem_1[840] = 64'd0;
	mem_1[841] = 64'd0;
	mem_1[842] = 64'd0;
	mem_1[843] = 64'd0;
	mem_1[844] = 64'd0;
	mem_1[845] = 64'd0;
	mem_1[846] = 64'd0;
	mem_1[847] = 64'd0;
	mem_1[848] = 64'd0;
	mem_1[849] = 64'd0;
	mem_1[850] = 64'd0;
	mem_1[851] = 64'd0;
	mem_1[852] = 64'd0;
	mem_1[853] = 64'd0;
	mem_1[854] = 64'd0;
	mem_1[855] = 64'd0;
	mem_1[856] = 64'd0;
	mem_1[857] = 64'd0;
	mem_1[858] = 64'd0;
	mem_1[859] = 64'd0;
	mem_1[860] = 64'd0;
	mem_1[861] = 64'd0;
	mem_1[862] = 64'd0;
	mem_1[863] = 64'd0;
	mem_1[864] = 64'd0;
	mem_1[865] = 64'd0;
	mem_1[866] = 64'd0;
	mem_1[867] = 64'd0;
	mem_1[868] = 64'd0;
	mem_1[869] = 64'd0;
	mem_1[870] = 64'd0;
	mem_1[871] = 64'd0;
	mem_1[872] = 64'd0;
	mem_1[873] = 64'd0;
	mem_1[874] = 64'd0;
	mem_1[875] = 64'd0;
	mem_1[876] = 64'd0;
	mem_1[877] = 64'd0;
	mem_1[878] = 64'd0;
	mem_1[879] = 64'd0;
	mem_1[880] = 64'd0;
	mem_1[881] = 64'd0;
	mem_1[882] = 64'd0;
	mem_1[883] = 64'd0;
	mem_1[884] = 64'd0;
	mem_1[885] = 64'd0;
	mem_1[886] = 64'd0;
	mem_1[887] = 64'd0;
	mem_1[888] = 64'd0;
	mem_1[889] = 64'd0;
	mem_1[890] = 64'd0;
	mem_1[891] = 64'd0;
	mem_1[892] = 64'd0;
	mem_1[893] = 64'd0;
	mem_1[894] = 64'd0;
	mem_1[895] = 64'd0;
	mem_1[896] = 64'd0;
	mem_1[897] = 64'd0;
	mem_1[898] = 64'd0;
	mem_1[899] = 64'd0;
	mem_1[900] = 64'd0;
	mem_1[901] = 64'd0;
	mem_1[902] = 64'd0;
	mem_1[903] = 64'd0;
	mem_1[904] = 64'd0;
	mem_1[905] = 64'd0;
	mem_1[906] = 64'd0;
	mem_1[907] = 64'd0;
	mem_1[908] = 64'd0;
	mem_1[909] = 64'd0;
	mem_1[910] = 64'd0;
	mem_1[911] = 64'd0;
	mem_1[912] = 64'd0;
	mem_1[913] = 64'd0;
	mem_1[914] = 64'd0;
	mem_1[915] = 64'd0;
	mem_1[916] = 64'd0;
	mem_1[917] = 64'd0;
	mem_1[918] = 64'd0;
	mem_1[919] = 64'd0;
	mem_1[920] = 64'd0;
	mem_1[921] = 64'd0;
	mem_1[922] = 64'd0;
	mem_1[923] = 64'd0;
	mem_1[924] = 64'd0;
	mem_1[925] = 64'd0;
	mem_1[926] = 64'd0;
	mem_1[927] = 64'd0;
	mem_1[928] = 64'd0;
	mem_1[929] = 64'd0;
	mem_1[930] = 64'd0;
	mem_1[931] = 64'd0;
	mem_1[932] = 64'd0;
	mem_1[933] = 64'd0;
	mem_1[934] = 64'd0;
	mem_1[935] = 64'd0;
	mem_1[936] = 64'd0;
	mem_1[937] = 64'd0;
	mem_1[938] = 64'd0;
	mem_1[939] = 64'd0;
	mem_1[940] = 64'd0;
	mem_1[941] = 64'd0;
	mem_1[942] = 64'd0;
	mem_1[943] = 64'd0;
	mem_1[944] = 64'd0;
	mem_1[945] = 64'd0;
	mem_1[946] = 64'd0;
	mem_1[947] = 64'd0;
	mem_1[948] = 64'd0;
	mem_1[949] = 64'd0;
	mem_1[950] = 64'd0;
	mem_1[951] = 64'd0;
	mem_1[952] = 64'd0;
	mem_1[953] = 64'd0;
	mem_1[954] = 64'd0;
	mem_1[955] = 64'd0;
	mem_1[956] = 64'd0;
	mem_1[957] = 64'd0;
	mem_1[958] = 64'd0;
	mem_1[959] = 64'd0;
	mem_1[960] = 64'd0;
	mem_1[961] = 64'd0;
	mem_1[962] = 64'd0;
	mem_1[963] = 64'd0;
	mem_1[964] = 64'd0;
	mem_1[965] = 64'd0;
	mem_1[966] = 64'd0;
	mem_1[967] = 64'd0;
	mem_1[968] = 64'd0;
	mem_1[969] = 64'd0;
	mem_1[970] = 64'd0;
	mem_1[971] = 64'd0;
	mem_1[972] = 64'd0;
	mem_1[973] = 64'd0;
	mem_1[974] = 64'd0;
	mem_1[975] = 64'd0;
	mem_1[976] = 64'd0;
	mem_1[977] = 64'd0;
	mem_1[978] = 64'd0;
	mem_1[979] = 64'd0;
	mem_1[980] = 64'd0;
	mem_1[981] = 64'd0;
	mem_1[982] = 64'd0;
	mem_1[983] = 64'd0;
	mem_1[984] = 64'd0;
	mem_1[985] = 64'd0;
	mem_1[986] = 64'd0;
	mem_1[987] = 64'd0;
	mem_1[988] = 64'd0;
	mem_1[989] = 64'd0;
	mem_1[990] = 64'd0;
	mem_1[991] = 64'd0;
	mem_1[992] = 64'd0;
	mem_1[993] = 64'd0;
	mem_1[994] = 64'd0;
	mem_1[995] = 64'd0;
	mem_1[996] = 64'd0;
	mem_1[997] = 64'd0;
	mem_1[998] = 64'd0;
	mem_1[999] = 64'd0;
	mem_1[1000] = 64'd0;
	mem_1[1001] = 64'd0;
	mem_1[1002] = 64'd0;
	mem_1[1003] = 64'd0;
	mem_1[1004] = 64'd0;
	mem_1[1005] = 64'd0;
	mem_1[1006] = 64'd0;
	mem_1[1007] = 64'd0;
	mem_1[1008] = 64'd0;
	mem_1[1009] = 64'd0;
	mem_1[1010] = 64'd0;
	mem_1[1011] = 64'd0;
	mem_1[1012] = 64'd0;
	mem_1[1013] = 64'd0;
	mem_1[1014] = 64'd0;
	mem_1[1015] = 64'd0;
	mem_1[1016] = 64'd0;
	mem_1[1017] = 64'd0;
	mem_1[1018] = 64'd0;
	mem_1[1019] = 64'd0;
	mem_1[1020] = 64'd0;
	mem_1[1021] = 64'd0;
	mem_1[1022] = 64'd0;
	mem_1[1023] = 64'd0;
	mem_2[0] = 64'd0;
	mem_2[1] = 64'd0;
	mem_2[2] = 64'd0;
	mem_2[3] = 64'd0;
	mem_2[4] = 64'd0;
	mem_2[5] = 64'd0;
	mem_2[6] = 64'd0;
	mem_2[7] = 64'd0;
	mem_2[8] = 64'd0;
	mem_2[9] = 64'd0;
	mem_2[10] = 64'd0;
	mem_2[11] = 64'd0;
	mem_2[12] = 64'd0;
	mem_2[13] = 64'd0;
	mem_2[14] = 64'd0;
	mem_2[15] = 64'd0;
	mem_2[16] = 64'd0;
	mem_2[17] = 64'd0;
	mem_2[18] = 64'd0;
	mem_2[19] = 64'd0;
	mem_2[20] = 64'd0;
	mem_2[21] = 64'd0;
	mem_2[22] = 64'd0;
	mem_2[23] = 64'd0;
	mem_2[24] = 64'd0;
	mem_2[25] = 64'd0;
	mem_2[26] = 64'd0;
	mem_2[27] = 64'd0;
	mem_2[28] = 64'd0;
	mem_2[29] = 64'd0;
	mem_2[30] = 64'd0;
	mem_2[31] = 64'd0;
	mem_2[32] = 64'd0;
	mem_2[33] = 64'd0;
	mem_2[34] = 64'd0;
	mem_2[35] = 64'd0;
	mem_2[36] = 64'd0;
	mem_2[37] = 64'd0;
	mem_2[38] = 64'd0;
	mem_2[39] = 64'd0;
	mem_2[40] = 64'd0;
	mem_2[41] = 64'd0;
	mem_2[42] = 64'd0;
	mem_2[43] = 64'd0;
	mem_2[44] = 64'd0;
	mem_2[45] = 64'd0;
	mem_2[46] = 64'd0;
	mem_2[47] = 64'd0;
	mem_2[48] = 64'd0;
	mem_2[49] = 64'd0;
	mem_2[50] = 64'd0;
	mem_2[51] = 64'd0;
	mem_2[52] = 64'd0;
	mem_2[53] = 64'd0;
	mem_2[54] = 64'd0;
	mem_2[55] = 64'd0;
	mem_2[56] = 64'd0;
	mem_2[57] = 64'd0;
	mem_2[58] = 64'd0;
	mem_2[59] = 64'd0;
	mem_2[60] = 64'd0;
	mem_2[61] = 64'd0;
	mem_2[62] = 64'd0;
	mem_2[63] = 64'd0;
	mem_2[64] = 64'd0;
	mem_2[65] = 64'd0;
	mem_2[66] = 64'd0;
	mem_2[67] = 64'd0;
	mem_2[68] = 64'd0;
	mem_2[69] = 64'd0;
	mem_2[70] = 64'd0;
	mem_2[71] = 64'd0;
	mem_2[72] = 64'd0;
	mem_2[73] = 64'd0;
	mem_2[74] = 64'd0;
	mem_2[75] = 64'd0;
	mem_2[76] = 64'd0;
	mem_2[77] = 64'd0;
	mem_2[78] = 64'd0;
	mem_2[79] = 64'd0;
	mem_2[80] = 64'd0;
	mem_2[81] = 64'd0;
	mem_2[82] = 64'd0;
	mem_2[83] = 64'd0;
	mem_2[84] = 64'd0;
	mem_2[85] = 64'd0;
	mem_2[86] = 64'd0;
	mem_2[87] = 64'd0;
	mem_2[88] = 64'd0;
	mem_2[89] = 64'd0;
	mem_2[90] = 64'd0;
	mem_2[91] = 64'd0;
	mem_2[92] = 64'd0;
	mem_2[93] = 64'd0;
	mem_2[94] = 64'd0;
	mem_2[95] = 64'd0;
	mem_2[96] = 64'd0;
	mem_2[97] = 64'd0;
	mem_2[98] = 64'd0;
	mem_2[99] = 64'd0;
	mem_2[100] = 64'd0;
	mem_2[101] = 64'd0;
	mem_2[102] = 64'd0;
	mem_2[103] = 64'd0;
	mem_2[104] = 64'd0;
	mem_2[105] = 64'd0;
	mem_2[106] = 64'd0;
	mem_2[107] = 64'd0;
	mem_2[108] = 64'd0;
	mem_2[109] = 64'd0;
	mem_2[110] = 64'd0;
	mem_2[111] = 64'd0;
	mem_2[112] = 64'd0;
	mem_2[113] = 64'd0;
	mem_2[114] = 64'd0;
	mem_2[115] = 64'd0;
	mem_2[116] = 64'd0;
	mem_2[117] = 64'd0;
	mem_2[118] = 64'd0;
	mem_2[119] = 64'd0;
	mem_2[120] = 64'd0;
	mem_2[121] = 64'd0;
	mem_2[122] = 64'd0;
	mem_2[123] = 64'd0;
	mem_2[124] = 64'd0;
	mem_2[125] = 64'd0;
	mem_2[126] = 64'd0;
	mem_2[127] = 64'd0;
	mem_2[128] = 64'd0;
	mem_2[129] = 64'd0;
	mem_2[130] = 64'd0;
	mem_2[131] = 64'd0;
	mem_2[132] = 64'd0;
	mem_2[133] = 64'd0;
	mem_2[134] = 64'd0;
	mem_2[135] = 64'd0;
	mem_2[136] = 64'd0;
	mem_2[137] = 64'd0;
	mem_2[138] = 64'd0;
	mem_2[139] = 64'd0;
	mem_2[140] = 64'd0;
	mem_2[141] = 64'd0;
	mem_2[142] = 64'd0;
	mem_2[143] = 64'd0;
	mem_2[144] = 64'd0;
	mem_2[145] = 64'd0;
	mem_2[146] = 64'd0;
	mem_2[147] = 64'd0;
	mem_2[148] = 64'd0;
	mem_2[149] = 64'd0;
	mem_2[150] = 64'd0;
	mem_2[151] = 64'd0;
	mem_2[152] = 64'd0;
	mem_2[153] = 64'd0;
	mem_2[154] = 64'd0;
	mem_2[155] = 64'd0;
	mem_2[156] = 64'd0;
	mem_2[157] = 64'd0;
	mem_2[158] = 64'd0;
	mem_2[159] = 64'd0;
	mem_2[160] = 64'd0;
	mem_2[161] = 64'd0;
	mem_2[162] = 64'd0;
	mem_2[163] = 64'd0;
	mem_2[164] = 64'd0;
	mem_2[165] = 64'd0;
	mem_2[166] = 64'd0;
	mem_2[167] = 64'd0;
	mem_2[168] = 64'd0;
	mem_2[169] = 64'd0;
	mem_2[170] = 64'd0;
	mem_2[171] = 64'd0;
	mem_2[172] = 64'd0;
	mem_2[173] = 64'd0;
	mem_2[174] = 64'd0;
	mem_2[175] = 64'd0;
	mem_2[176] = 64'd0;
	mem_2[177] = 64'd0;
	mem_2[178] = 64'd0;
	mem_2[179] = 64'd0;
	mem_2[180] = 64'd0;
	mem_2[181] = 64'd0;
	mem_2[182] = 64'd0;
	mem_2[183] = 64'd0;
	mem_2[184] = 64'd0;
	mem_2[185] = 64'd0;
	mem_2[186] = 64'd0;
	mem_2[187] = 64'd0;
	mem_2[188] = 64'd0;
	mem_2[189] = 64'd0;
	mem_2[190] = 64'd0;
	mem_2[191] = 64'd0;
	mem_2[192] = 64'd0;
	mem_2[193] = 64'd0;
	mem_2[194] = 64'd0;
	mem_2[195] = 64'd0;
	mem_2[196] = 64'd0;
	mem_2[197] = 64'd0;
	mem_2[198] = 64'd0;
	mem_2[199] = 64'd0;
	mem_2[200] = 64'd0;
	mem_2[201] = 64'd0;
	mem_2[202] = 64'd0;
	mem_2[203] = 64'd0;
	mem_2[204] = 64'd0;
	mem_2[205] = 64'd0;
	mem_2[206] = 64'd0;
	mem_2[207] = 64'd0;
	mem_2[208] = 64'd0;
	mem_2[209] = 64'd0;
	mem_2[210] = 64'd0;
	mem_2[211] = 64'd0;
	mem_2[212] = 64'd0;
	mem_2[213] = 64'd0;
	mem_2[214] = 64'd0;
	mem_2[215] = 64'd0;
	mem_2[216] = 64'd0;
	mem_2[217] = 64'd0;
	mem_2[218] = 64'd0;
	mem_2[219] = 64'd0;
	mem_2[220] = 64'd0;
	mem_2[221] = 64'd0;
	mem_2[222] = 64'd0;
	mem_2[223] = 64'd0;
	mem_2[224] = 64'd0;
	mem_2[225] = 64'd0;
	mem_2[226] = 64'd0;
	mem_2[227] = 64'd0;
	mem_2[228] = 64'd0;
	mem_2[229] = 64'd0;
	mem_2[230] = 64'd0;
	mem_2[231] = 64'd0;
	mem_2[232] = 64'd0;
	mem_2[233] = 64'd0;
	mem_2[234] = 64'd0;
	mem_2[235] = 64'd0;
	mem_2[236] = 64'd0;
	mem_2[237] = 64'd0;
	mem_2[238] = 64'd0;
	mem_2[239] = 64'd0;
	mem_2[240] = 64'd0;
	mem_2[241] = 64'd0;
	mem_2[242] = 64'd0;
	mem_2[243] = 64'd0;
	mem_2[244] = 64'd0;
	mem_2[245] = 64'd0;
	mem_2[246] = 64'd0;
	mem_2[247] = 64'd0;
	mem_2[248] = 64'd0;
	mem_2[249] = 64'd0;
	mem_2[250] = 64'd0;
	mem_2[251] = 64'd0;
	mem_2[252] = 64'd0;
	mem_2[253] = 64'd0;
	mem_2[254] = 64'd0;
	mem_2[255] = 64'd0;
	mem_2[256] = 64'd0;
	mem_2[257] = 64'd0;
	mem_2[258] = 64'd0;
	mem_2[259] = 64'd0;
	mem_2[260] = 64'd0;
	mem_2[261] = 64'd0;
	mem_2[262] = 64'd0;
	mem_2[263] = 64'd0;
	mem_2[264] = 64'd0;
	mem_2[265] = 64'd0;
	mem_2[266] = 64'd0;
	mem_2[267] = 64'd0;
	mem_2[268] = 64'd0;
	mem_2[269] = 64'd0;
	mem_2[270] = 64'd0;
	mem_2[271] = 64'd0;
	mem_2[272] = 64'd0;
	mem_2[273] = 64'd0;
	mem_2[274] = 64'd0;
	mem_2[275] = 64'd0;
	mem_2[276] = 64'd0;
	mem_2[277] = 64'd0;
	mem_2[278] = 64'd0;
	mem_2[279] = 64'd0;
	mem_2[280] = 64'd0;
	mem_2[281] = 64'd0;
	mem_2[282] = 64'd0;
	mem_2[283] = 64'd0;
	mem_2[284] = 64'd0;
	mem_2[285] = 64'd0;
	mem_2[286] = 64'd0;
	mem_2[287] = 64'd0;
	mem_2[288] = 64'd0;
	mem_2[289] = 64'd0;
	mem_2[290] = 64'd0;
	mem_2[291] = 64'd0;
	mem_2[292] = 64'd0;
	mem_2[293] = 64'd0;
	mem_2[294] = 64'd0;
	mem_2[295] = 64'd0;
	mem_2[296] = 64'd0;
	mem_2[297] = 64'd0;
	mem_2[298] = 64'd0;
	mem_2[299] = 64'd0;
	mem_2[300] = 64'd0;
	mem_2[301] = 64'd0;
	mem_2[302] = 64'd0;
	mem_2[303] = 64'd0;
	mem_2[304] = 64'd0;
	mem_2[305] = 64'd0;
	mem_2[306] = 64'd0;
	mem_2[307] = 64'd0;
	mem_2[308] = 64'd0;
	mem_2[309] = 64'd0;
	mem_2[310] = 64'd0;
	mem_2[311] = 64'd0;
	mem_2[312] = 64'd0;
	mem_2[313] = 64'd0;
	mem_2[314] = 64'd0;
	mem_2[315] = 64'd0;
	mem_2[316] = 64'd0;
	mem_2[317] = 64'd0;
	mem_2[318] = 64'd0;
	mem_2[319] = 64'd0;
	mem_2[320] = 64'd0;
	mem_2[321] = 64'd0;
	mem_2[322] = 64'd0;
	mem_2[323] = 64'd0;
	mem_2[324] = 64'd0;
	mem_2[325] = 64'd0;
	mem_2[326] = 64'd0;
	mem_2[327] = 64'd0;
	mem_2[328] = 64'd0;
	mem_2[329] = 64'd0;
	mem_2[330] = 64'd0;
	mem_2[331] = 64'd0;
	mem_2[332] = 64'd0;
	mem_2[333] = 64'd0;
	mem_2[334] = 64'd0;
	mem_2[335] = 64'd0;
	mem_2[336] = 64'd0;
	mem_2[337] = 64'd0;
	mem_2[338] = 64'd0;
	mem_2[339] = 64'd0;
	mem_2[340] = 64'd0;
	mem_2[341] = 64'd0;
	mem_2[342] = 64'd0;
	mem_2[343] = 64'd0;
	mem_2[344] = 64'd0;
	mem_2[345] = 64'd0;
	mem_2[346] = 64'd0;
	mem_2[347] = 64'd0;
	mem_2[348] = 64'd0;
	mem_2[349] = 64'd0;
	mem_2[350] = 64'd0;
	mem_2[351] = 64'd0;
	mem_2[352] = 64'd0;
	mem_2[353] = 64'd0;
	mem_2[354] = 64'd0;
	mem_2[355] = 64'd0;
	mem_2[356] = 64'd0;
	mem_2[357] = 64'd0;
	mem_2[358] = 64'd0;
	mem_2[359] = 64'd0;
	mem_2[360] = 64'd0;
	mem_2[361] = 64'd0;
	mem_2[362] = 64'd0;
	mem_2[363] = 64'd0;
	mem_2[364] = 64'd0;
	mem_2[365] = 64'd0;
	mem_2[366] = 64'd0;
	mem_2[367] = 64'd0;
	mem_2[368] = 64'd0;
	mem_2[369] = 64'd0;
	mem_2[370] = 64'd0;
	mem_2[371] = 64'd0;
	mem_2[372] = 64'd0;
	mem_2[373] = 64'd0;
	mem_2[374] = 64'd0;
	mem_2[375] = 64'd0;
	mem_2[376] = 64'd0;
	mem_2[377] = 64'd0;
	mem_2[378] = 64'd0;
	mem_2[379] = 64'd0;
	mem_2[380] = 64'd0;
	mem_2[381] = 64'd0;
	mem_2[382] = 64'd0;
	mem_2[383] = 64'd0;
	mem_2[384] = 64'd0;
	mem_2[385] = 64'd0;
	mem_2[386] = 64'd0;
	mem_2[387] = 64'd0;
	mem_2[388] = 64'd0;
	mem_2[389] = 64'd0;
	mem_2[390] = 64'd0;
	mem_2[391] = 64'd0;
	mem_2[392] = 64'd0;
	mem_2[393] = 64'd0;
	mem_2[394] = 64'd0;
	mem_2[395] = 64'd0;
	mem_2[396] = 64'd0;
	mem_2[397] = 64'd0;
	mem_2[398] = 64'd0;
	mem_2[399] = 64'd0;
	mem_2[400] = 64'd0;
	mem_2[401] = 64'd0;
	mem_2[402] = 64'd0;
	mem_2[403] = 64'd0;
	mem_2[404] = 64'd0;
	mem_2[405] = 64'd0;
	mem_2[406] = 64'd0;
	mem_2[407] = 64'd0;
	mem_2[408] = 64'd0;
	mem_2[409] = 64'd0;
	mem_2[410] = 64'd0;
	mem_2[411] = 64'd0;
	mem_2[412] = 64'd0;
	mem_2[413] = 64'd0;
	mem_2[414] = 64'd0;
	mem_2[415] = 64'd0;
	mem_2[416] = 64'd0;
	mem_2[417] = 64'd0;
	mem_2[418] = 64'd0;
	mem_2[419] = 64'd0;
	mem_2[420] = 64'd0;
	mem_2[421] = 64'd0;
	mem_2[422] = 64'd0;
	mem_2[423] = 64'd0;
	mem_2[424] = 64'd0;
	mem_2[425] = 64'd0;
	mem_2[426] = 64'd0;
	mem_2[427] = 64'd0;
	mem_2[428] = 64'd0;
	mem_2[429] = 64'd0;
	mem_2[430] = 64'd0;
	mem_2[431] = 64'd0;
	mem_2[432] = 64'd0;
	mem_2[433] = 64'd0;
	mem_2[434] = 64'd0;
	mem_2[435] = 64'd0;
	mem_2[436] = 64'd0;
	mem_2[437] = 64'd0;
	mem_2[438] = 64'd0;
	mem_2[439] = 64'd0;
	mem_2[440] = 64'd0;
	mem_2[441] = 64'd0;
	mem_2[442] = 64'd0;
	mem_2[443] = 64'd0;
	mem_2[444] = 64'd0;
	mem_2[445] = 64'd0;
	mem_2[446] = 64'd0;
	mem_2[447] = 64'd0;
	mem_2[448] = 64'd0;
	mem_2[449] = 64'd0;
	mem_2[450] = 64'd0;
	mem_2[451] = 64'd0;
	mem_2[452] = 64'd0;
	mem_2[453] = 64'd0;
	mem_2[454] = 64'd0;
	mem_2[455] = 64'd0;
	mem_2[456] = 64'd0;
	mem_2[457] = 64'd0;
	mem_2[458] = 64'd0;
	mem_2[459] = 64'd0;
	mem_2[460] = 64'd0;
	mem_2[461] = 64'd0;
	mem_2[462] = 64'd0;
	mem_2[463] = 64'd0;
	mem_2[464] = 64'd0;
	mem_2[465] = 64'd0;
	mem_2[466] = 64'd0;
	mem_2[467] = 64'd0;
	mem_2[468] = 64'd0;
	mem_2[469] = 64'd0;
	mem_2[470] = 64'd0;
	mem_2[471] = 64'd0;
	mem_2[472] = 64'd0;
	mem_2[473] = 64'd0;
	mem_2[474] = 64'd0;
	mem_2[475] = 64'd0;
	mem_2[476] = 64'd0;
	mem_2[477] = 64'd0;
	mem_2[478] = 64'd0;
	mem_2[479] = 64'd0;
	mem_2[480] = 64'd0;
	mem_2[481] = 64'd0;
	mem_2[482] = 64'd0;
	mem_2[483] = 64'd0;
	mem_2[484] = 64'd0;
	mem_2[485] = 64'd0;
	mem_2[486] = 64'd0;
	mem_2[487] = 64'd0;
	mem_2[488] = 64'd0;
	mem_2[489] = 64'd0;
	mem_2[490] = 64'd0;
	mem_2[491] = 64'd0;
	mem_2[492] = 64'd0;
	mem_2[493] = 64'd0;
	mem_2[494] = 64'd0;
	mem_2[495] = 64'd0;
	mem_2[496] = 64'd0;
	mem_2[497] = 64'd0;
	mem_2[498] = 64'd0;
	mem_2[499] = 64'd0;
	mem_2[500] = 64'd0;
	mem_2[501] = 64'd0;
	mem_2[502] = 64'd0;
	mem_2[503] = 64'd0;
	mem_2[504] = 64'd0;
	mem_2[505] = 64'd0;
	mem_2[506] = 64'd0;
	mem_2[507] = 64'd0;
	mem_2[508] = 64'd0;
	mem_2[509] = 64'd0;
	mem_2[510] = 64'd0;
	mem_2[511] = 64'd0;
	mem_2[512] = 64'd0;
	mem_2[513] = 64'd0;
	mem_2[514] = 64'd0;
	mem_2[515] = 64'd0;
	mem_2[516] = 64'd0;
	mem_2[517] = 64'd0;
	mem_2[518] = 64'd0;
	mem_2[519] = 64'd0;
	mem_2[520] = 64'd0;
	mem_2[521] = 64'd0;
	mem_2[522] = 64'd0;
	mem_2[523] = 64'd0;
	mem_2[524] = 64'd0;
	mem_2[525] = 64'd0;
	mem_2[526] = 64'd0;
	mem_2[527] = 64'd0;
	mem_2[528] = 64'd0;
	mem_2[529] = 64'd0;
	mem_2[530] = 64'd0;
	mem_2[531] = 64'd0;
	mem_2[532] = 64'd0;
	mem_2[533] = 64'd0;
	mem_2[534] = 64'd0;
	mem_2[535] = 64'd0;
	mem_2[536] = 64'd0;
	mem_2[537] = 64'd0;
	mem_2[538] = 64'd0;
	mem_2[539] = 64'd0;
	mem_2[540] = 64'd0;
	mem_2[541] = 64'd0;
	mem_2[542] = 64'd0;
	mem_2[543] = 64'd0;
	mem_2[544] = 64'd0;
	mem_2[545] = 64'd0;
	mem_2[546] = 64'd0;
	mem_2[547] = 64'd0;
	mem_2[548] = 64'd0;
	mem_2[549] = 64'd0;
	mem_2[550] = 64'd0;
	mem_2[551] = 64'd0;
	mem_2[552] = 64'd0;
	mem_2[553] = 64'd0;
	mem_2[554] = 64'd0;
	mem_2[555] = 64'd0;
	mem_2[556] = 64'd0;
	mem_2[557] = 64'd0;
	mem_2[558] = 64'd0;
	mem_2[559] = 64'd0;
	mem_2[560] = 64'd0;
	mem_2[561] = 64'd0;
	mem_2[562] = 64'd0;
	mem_2[563] = 64'd0;
	mem_2[564] = 64'd0;
	mem_2[565] = 64'd0;
	mem_2[566] = 64'd0;
	mem_2[567] = 64'd0;
	mem_2[568] = 64'd0;
	mem_2[569] = 64'd0;
	mem_2[570] = 64'd0;
	mem_2[571] = 64'd0;
	mem_2[572] = 64'd0;
	mem_2[573] = 64'd0;
	mem_2[574] = 64'd0;
	mem_2[575] = 64'd0;
	mem_2[576] = 64'd0;
	mem_2[577] = 64'd0;
	mem_2[578] = 64'd0;
	mem_2[579] = 64'd0;
	mem_2[580] = 64'd0;
	mem_2[581] = 64'd0;
	mem_2[582] = 64'd0;
	mem_2[583] = 64'd0;
	mem_2[584] = 64'd0;
	mem_2[585] = 64'd0;
	mem_2[586] = 64'd0;
	mem_2[587] = 64'd0;
	mem_2[588] = 64'd0;
	mem_2[589] = 64'd0;
	mem_2[590] = 64'd0;
	mem_2[591] = 64'd0;
	mem_2[592] = 64'd0;
	mem_2[593] = 64'd0;
	mem_2[594] = 64'd0;
	mem_2[595] = 64'd0;
	mem_2[596] = 64'd0;
	mem_2[597] = 64'd0;
	mem_2[598] = 64'd0;
	mem_2[599] = 64'd0;
	mem_2[600] = 64'd0;
	mem_2[601] = 64'd0;
	mem_2[602] = 64'd0;
	mem_2[603] = 64'd0;
	mem_2[604] = 64'd0;
	mem_2[605] = 64'd0;
	mem_2[606] = 64'd0;
	mem_2[607] = 64'd0;
	mem_2[608] = 64'd0;
	mem_2[609] = 64'd0;
	mem_2[610] = 64'd0;
	mem_2[611] = 64'd0;
	mem_2[612] = 64'd0;
	mem_2[613] = 64'd0;
	mem_2[614] = 64'd0;
	mem_2[615] = 64'd0;
	mem_2[616] = 64'd0;
	mem_2[617] = 64'd0;
	mem_2[618] = 64'd0;
	mem_2[619] = 64'd0;
	mem_2[620] = 64'd0;
	mem_2[621] = 64'd0;
	mem_2[622] = 64'd0;
	mem_2[623] = 64'd0;
	mem_2[624] = 64'd0;
	mem_2[625] = 64'd0;
	mem_2[626] = 64'd0;
	mem_2[627] = 64'd0;
	mem_2[628] = 64'd0;
	mem_2[629] = 64'd0;
	mem_2[630] = 64'd0;
	mem_2[631] = 64'd0;
	mem_2[632] = 64'd0;
	mem_2[633] = 64'd0;
	mem_2[634] = 64'd0;
	mem_2[635] = 64'd0;
	mem_2[636] = 64'd0;
	mem_2[637] = 64'd0;
	mem_2[638] = 64'd0;
	mem_2[639] = 64'd0;
	mem_2[640] = 64'd0;
	mem_2[641] = 64'd0;
	mem_2[642] = 64'd0;
	mem_2[643] = 64'd0;
	mem_2[644] = 64'd0;
	mem_2[645] = 64'd0;
	mem_2[646] = 64'd0;
	mem_2[647] = 64'd0;
	mem_2[648] = 64'd0;
	mem_2[649] = 64'd0;
	mem_2[650] = 64'd0;
	mem_2[651] = 64'd0;
	mem_2[652] = 64'd0;
	mem_2[653] = 64'd0;
	mem_2[654] = 64'd0;
	mem_2[655] = 64'd0;
	mem_2[656] = 64'd0;
	mem_2[657] = 64'd0;
	mem_2[658] = 64'd0;
	mem_2[659] = 64'd0;
	mem_2[660] = 64'd0;
	mem_2[661] = 64'd0;
	mem_2[662] = 64'd0;
	mem_2[663] = 64'd0;
	mem_2[664] = 64'd0;
	mem_2[665] = 64'd0;
	mem_2[666] = 64'd0;
	mem_2[667] = 64'd0;
	mem_2[668] = 64'd0;
	mem_2[669] = 64'd0;
	mem_2[670] = 64'd0;
	mem_2[671] = 64'd0;
	mem_2[672] = 64'd0;
	mem_2[673] = 64'd0;
	mem_2[674] = 64'd0;
	mem_2[675] = 64'd0;
	mem_2[676] = 64'd0;
	mem_2[677] = 64'd0;
	mem_2[678] = 64'd0;
	mem_2[679] = 64'd0;
	mem_2[680] = 64'd0;
	mem_2[681] = 64'd0;
	mem_2[682] = 64'd0;
	mem_2[683] = 64'd0;
	mem_2[684] = 64'd0;
	mem_2[685] = 64'd0;
	mem_2[686] = 64'd0;
	mem_2[687] = 64'd0;
	mem_2[688] = 64'd0;
	mem_2[689] = 64'd0;
	mem_2[690] = 64'd0;
	mem_2[691] = 64'd0;
	mem_2[692] = 64'd0;
	mem_2[693] = 64'd0;
	mem_2[694] = 64'd0;
	mem_2[695] = 64'd0;
	mem_2[696] = 64'd0;
	mem_2[697] = 64'd0;
	mem_2[698] = 64'd0;
	mem_2[699] = 64'd0;
	mem_2[700] = 64'd0;
	mem_2[701] = 64'd0;
	mem_2[702] = 64'd0;
	mem_2[703] = 64'd0;
	mem_2[704] = 64'd0;
	mem_2[705] = 64'd0;
	mem_2[706] = 64'd0;
	mem_2[707] = 64'd0;
	mem_2[708] = 64'd0;
	mem_2[709] = 64'd0;
	mem_2[710] = 64'd0;
	mem_2[711] = 64'd0;
	mem_2[712] = 64'd0;
	mem_2[713] = 64'd0;
	mem_2[714] = 64'd0;
	mem_2[715] = 64'd0;
	mem_2[716] = 64'd0;
	mem_2[717] = 64'd0;
	mem_2[718] = 64'd0;
	mem_2[719] = 64'd0;
	mem_2[720] = 64'd0;
	mem_2[721] = 64'd0;
	mem_2[722] = 64'd0;
	mem_2[723] = 64'd0;
	mem_2[724] = 64'd0;
	mem_2[725] = 64'd0;
	mem_2[726] = 64'd0;
	mem_2[727] = 64'd0;
	mem_2[728] = 64'd0;
	mem_2[729] = 64'd0;
	mem_2[730] = 64'd0;
	mem_2[731] = 64'd0;
	mem_2[732] = 64'd0;
	mem_2[733] = 64'd0;
	mem_2[734] = 64'd0;
	mem_2[735] = 64'd0;
	mem_2[736] = 64'd0;
	mem_2[737] = 64'd0;
	mem_2[738] = 64'd0;
	mem_2[739] = 64'd0;
	mem_2[740] = 64'd0;
	mem_2[741] = 64'd0;
	mem_2[742] = 64'd0;
	mem_2[743] = 64'd0;
	mem_2[744] = 64'd0;
	mem_2[745] = 64'd0;
	mem_2[746] = 64'd0;
	mem_2[747] = 64'd0;
	mem_2[748] = 64'd0;
	mem_2[749] = 64'd0;
	mem_2[750] = 64'd0;
	mem_2[751] = 64'd0;
	mem_2[752] = 64'd0;
	mem_2[753] = 64'd0;
	mem_2[754] = 64'd0;
	mem_2[755] = 64'd0;
	mem_2[756] = 64'd0;
	mem_2[757] = 64'd0;
	mem_2[758] = 64'd0;
	mem_2[759] = 64'd0;
	mem_2[760] = 64'd0;
	mem_2[761] = 64'd0;
	mem_2[762] = 64'd0;
	mem_2[763] = 64'd0;
	mem_2[764] = 64'd0;
	mem_2[765] = 64'd0;
	mem_2[766] = 64'd0;
	mem_2[767] = 64'd0;
	mem_2[768] = 64'd0;
	mem_2[769] = 64'd0;
	mem_2[770] = 64'd0;
	mem_2[771] = 64'd0;
	mem_2[772] = 64'd0;
	mem_2[773] = 64'd0;
	mem_2[774] = 64'd0;
	mem_2[775] = 64'd0;
	mem_2[776] = 64'd0;
	mem_2[777] = 64'd0;
	mem_2[778] = 64'd0;
	mem_2[779] = 64'd0;
	mem_2[780] = 64'd0;
	mem_2[781] = 64'd0;
	mem_2[782] = 64'd0;
	mem_2[783] = 64'd0;
	mem_2[784] = 64'd0;
	mem_2[785] = 64'd0;
	mem_2[786] = 64'd0;
	mem_2[787] = 64'd0;
	mem_2[788] = 64'd0;
	mem_2[789] = 64'd0;
	mem_2[790] = 64'd0;
	mem_2[791] = 64'd0;
	mem_2[792] = 64'd0;
	mem_2[793] = 64'd0;
	mem_2[794] = 64'd0;
	mem_2[795] = 64'd0;
	mem_2[796] = 64'd0;
	mem_2[797] = 64'd0;
	mem_2[798] = 64'd0;
	mem_2[799] = 64'd0;
	mem_2[800] = 64'd0;
	mem_2[801] = 64'd0;
	mem_2[802] = 64'd0;
	mem_2[803] = 64'd0;
	mem_2[804] = 64'd0;
	mem_2[805] = 64'd0;
	mem_2[806] = 64'd0;
	mem_2[807] = 64'd0;
	mem_2[808] = 64'd0;
	mem_2[809] = 64'd0;
	mem_2[810] = 64'd0;
	mem_2[811] = 64'd0;
	mem_2[812] = 64'd0;
	mem_2[813] = 64'd0;
	mem_2[814] = 64'd0;
	mem_2[815] = 64'd0;
	mem_2[816] = 64'd0;
	mem_2[817] = 64'd0;
	mem_2[818] = 64'd0;
	mem_2[819] = 64'd0;
	mem_2[820] = 64'd0;
	mem_2[821] = 64'd0;
	mem_2[822] = 64'd0;
	mem_2[823] = 64'd0;
	mem_2[824] = 64'd0;
	mem_2[825] = 64'd0;
	mem_2[826] = 64'd0;
	mem_2[827] = 64'd0;
	mem_2[828] = 64'd0;
	mem_2[829] = 64'd0;
	mem_2[830] = 64'd0;
	mem_2[831] = 64'd0;
	mem_2[832] = 64'd0;
	mem_2[833] = 64'd0;
	mem_2[834] = 64'd0;
	mem_2[835] = 64'd0;
	mem_2[836] = 64'd0;
	mem_2[837] = 64'd0;
	mem_2[838] = 64'd0;
	mem_2[839] = 64'd0;
	mem_2[840] = 64'd0;
	mem_2[841] = 64'd0;
	mem_2[842] = 64'd0;
	mem_2[843] = 64'd0;
	mem_2[844] = 64'd0;
	mem_2[845] = 64'd0;
	mem_2[846] = 64'd0;
	mem_2[847] = 64'd0;
	mem_2[848] = 64'd0;
	mem_2[849] = 64'd0;
	mem_2[850] = 64'd0;
	mem_2[851] = 64'd0;
	mem_2[852] = 64'd0;
	mem_2[853] = 64'd0;
	mem_2[854] = 64'd0;
	mem_2[855] = 64'd0;
	mem_2[856] = 64'd0;
	mem_2[857] = 64'd0;
	mem_2[858] = 64'd0;
	mem_2[859] = 64'd0;
	mem_2[860] = 64'd0;
	mem_2[861] = 64'd0;
	mem_2[862] = 64'd0;
	mem_2[863] = 64'd0;
	mem_2[864] = 64'd0;
	mem_2[865] = 64'd0;
	mem_2[866] = 64'd0;
	mem_2[867] = 64'd0;
	mem_2[868] = 64'd0;
	mem_2[869] = 64'd0;
	mem_2[870] = 64'd0;
	mem_2[871] = 64'd0;
	mem_2[872] = 64'd0;
	mem_2[873] = 64'd0;
	mem_2[874] = 64'd0;
	mem_2[875] = 64'd0;
	mem_2[876] = 64'd0;
	mem_2[877] = 64'd0;
	mem_2[878] = 64'd0;
	mem_2[879] = 64'd0;
	mem_2[880] = 64'd0;
	mem_2[881] = 64'd0;
	mem_2[882] = 64'd0;
	mem_2[883] = 64'd0;
	mem_2[884] = 64'd0;
	mem_2[885] = 64'd0;
	mem_2[886] = 64'd0;
	mem_2[887] = 64'd0;
	mem_2[888] = 64'd0;
	mem_2[889] = 64'd0;
	mem_2[890] = 64'd0;
	mem_2[891] = 64'd0;
	mem_2[892] = 64'd0;
	mem_2[893] = 64'd0;
	mem_2[894] = 64'd0;
	mem_2[895] = 64'd0;
	mem_2[896] = 64'd0;
	mem_2[897] = 64'd0;
	mem_2[898] = 64'd0;
	mem_2[899] = 64'd0;
	mem_2[900] = 64'd0;
	mem_2[901] = 64'd0;
	mem_2[902] = 64'd0;
	mem_2[903] = 64'd0;
	mem_2[904] = 64'd0;
	mem_2[905] = 64'd0;
	mem_2[906] = 64'd0;
	mem_2[907] = 64'd0;
	mem_2[908] = 64'd0;
	mem_2[909] = 64'd0;
	mem_2[910] = 64'd0;
	mem_2[911] = 64'd0;
	mem_2[912] = 64'd0;
	mem_2[913] = 64'd0;
	mem_2[914] = 64'd0;
	mem_2[915] = 64'd0;
	mem_2[916] = 64'd0;
	mem_2[917] = 64'd0;
	mem_2[918] = 64'd0;
	mem_2[919] = 64'd0;
	mem_2[920] = 64'd0;
	mem_2[921] = 64'd0;
	mem_2[922] = 64'd0;
	mem_2[923] = 64'd0;
	mem_2[924] = 64'd0;
	mem_2[925] = 64'd0;
	mem_2[926] = 64'd0;
	mem_2[927] = 64'd0;
	mem_2[928] = 64'd0;
	mem_2[929] = 64'd0;
	mem_2[930] = 64'd0;
	mem_2[931] = 64'd0;
	mem_2[932] = 64'd0;
	mem_2[933] = 64'd0;
	mem_2[934] = 64'd0;
	mem_2[935] = 64'd0;
	mem_2[936] = 64'd0;
	mem_2[937] = 64'd0;
	mem_2[938] = 64'd0;
	mem_2[939] = 64'd0;
	mem_2[940] = 64'd0;
	mem_2[941] = 64'd0;
	mem_2[942] = 64'd0;
	mem_2[943] = 64'd0;
	mem_2[944] = 64'd0;
	mem_2[945] = 64'd0;
	mem_2[946] = 64'd0;
	mem_2[947] = 64'd0;
	mem_2[948] = 64'd0;
	mem_2[949] = 64'd0;
	mem_2[950] = 64'd0;
	mem_2[951] = 64'd0;
	mem_2[952] = 64'd0;
	mem_2[953] = 64'd0;
	mem_2[954] = 64'd0;
	mem_2[955] = 64'd0;
	mem_2[956] = 64'd0;
	mem_2[957] = 64'd0;
	mem_2[958] = 64'd0;
	mem_2[959] = 64'd0;
	mem_2[960] = 64'd0;
	mem_2[961] = 64'd0;
	mem_2[962] = 64'd0;
	mem_2[963] = 64'd0;
	mem_2[964] = 64'd0;
	mem_2[965] = 64'd0;
	mem_2[966] = 64'd0;
	mem_2[967] = 64'd0;
	mem_2[968] = 64'd0;
	mem_2[969] = 64'd0;
	mem_2[970] = 64'd0;
	mem_2[971] = 64'd0;
	mem_2[972] = 64'd0;
	mem_2[973] = 64'd0;
	mem_2[974] = 64'd0;
	mem_2[975] = 64'd0;
	mem_2[976] = 64'd0;
	mem_2[977] = 64'd0;
	mem_2[978] = 64'd0;
	mem_2[979] = 64'd0;
	mem_2[980] = 64'd0;
	mem_2[981] = 64'd0;
	mem_2[982] = 64'd0;
	mem_2[983] = 64'd0;
	mem_2[984] = 64'd0;
	mem_2[985] = 64'd0;
	mem_2[986] = 64'd0;
	mem_2[987] = 64'd0;
	mem_2[988] = 64'd0;
	mem_2[989] = 64'd0;
	mem_2[990] = 64'd0;
	mem_2[991] = 64'd0;
	mem_2[992] = 64'd0;
	mem_2[993] = 64'd0;
	mem_2[994] = 64'd0;
	mem_2[995] = 64'd0;
	mem_2[996] = 64'd0;
	mem_2[997] = 64'd0;
	mem_2[998] = 64'd0;
	mem_2[999] = 64'd0;
	mem_2[1000] = 64'd0;
	mem_2[1001] = 64'd0;
	mem_2[1002] = 64'd0;
	mem_2[1003] = 64'd0;
	mem_2[1004] = 64'd0;
	mem_2[1005] = 64'd0;
	mem_2[1006] = 64'd0;
	mem_2[1007] = 64'd0;
	mem_2[1008] = 64'd0;
	mem_2[1009] = 64'd0;
	mem_2[1010] = 64'd0;
	mem_2[1011] = 64'd0;
	mem_2[1012] = 64'd0;
	mem_2[1013] = 64'd0;
	mem_2[1014] = 64'd0;
	mem_2[1015] = 64'd0;
	mem_2[1016] = 64'd0;
	mem_2[1017] = 64'd0;
	mem_2[1018] = 64'd0;
	mem_2[1019] = 64'd0;
	mem_2[1020] = 64'd0;
	mem_2[1021] = 64'd0;
	mem_2[1022] = 64'd0;
	mem_2[1023] = 64'd0;
	mem_3[0] = 64'd0;
	mem_3[1] = 64'd0;
	mem_3[2] = 64'd0;
	mem_3[3] = 64'd0;
	mem_3[4] = 64'd0;
	mem_3[5] = 64'd0;
	mem_3[6] = 64'd0;
	mem_3[7] = 64'd0;
	mem_3[8] = 64'd0;
	mem_3[9] = 64'd0;
	mem_3[10] = 64'd0;
	mem_3[11] = 64'd0;
	mem_3[12] = 64'd0;
	mem_3[13] = 64'd0;
	mem_3[14] = 64'd0;
	mem_3[15] = 64'd0;
	mem_3[16] = 64'd0;
	mem_3[17] = 64'd0;
	mem_3[18] = 64'd0;
	mem_3[19] = 64'd0;
	mem_3[20] = 64'd0;
	mem_3[21] = 64'd0;
	mem_3[22] = 64'd0;
	mem_3[23] = 64'd0;
	mem_3[24] = 64'd0;
	mem_3[25] = 64'd0;
	mem_3[26] = 64'd0;
	mem_3[27] = 64'd0;
	mem_3[28] = 64'd0;
	mem_3[29] = 64'd0;
	mem_3[30] = 64'd0;
	mem_3[31] = 64'd0;
	mem_3[32] = 64'd0;
	mem_3[33] = 64'd0;
	mem_3[34] = 64'd0;
	mem_3[35] = 64'd0;
	mem_3[36] = 64'd0;
	mem_3[37] = 64'd0;
	mem_3[38] = 64'd0;
	mem_3[39] = 64'd0;
	mem_3[40] = 64'd0;
	mem_3[41] = 64'd0;
	mem_3[42] = 64'd0;
	mem_3[43] = 64'd0;
	mem_3[44] = 64'd0;
	mem_3[45] = 64'd0;
	mem_3[46] = 64'd0;
	mem_3[47] = 64'd0;
	mem_3[48] = 64'd0;
	mem_3[49] = 64'd0;
	mem_3[50] = 64'd0;
	mem_3[51] = 64'd0;
	mem_3[52] = 64'd0;
	mem_3[53] = 64'd0;
	mem_3[54] = 64'd0;
	mem_3[55] = 64'd0;
	mem_3[56] = 64'd0;
	mem_3[57] = 64'd0;
	mem_3[58] = 64'd0;
	mem_3[59] = 64'd0;
	mem_3[60] = 64'd0;
	mem_3[61] = 64'd0;
	mem_3[62] = 64'd0;
	mem_3[63] = 64'd0;
	mem_3[64] = 64'd0;
	mem_3[65] = 64'd0;
	mem_3[66] = 64'd0;
	mem_3[67] = 64'd0;
	mem_3[68] = 64'd0;
	mem_3[69] = 64'd0;
	mem_3[70] = 64'd0;
	mem_3[71] = 64'd0;
	mem_3[72] = 64'd0;
	mem_3[73] = 64'd0;
	mem_3[74] = 64'd0;
	mem_3[75] = 64'd0;
	mem_3[76] = 64'd0;
	mem_3[77] = 64'd0;
	mem_3[78] = 64'd0;
	mem_3[79] = 64'd0;
	mem_3[80] = 64'd0;
	mem_3[81] = 64'd0;
	mem_3[82] = 64'd0;
	mem_3[83] = 64'd0;
	mem_3[84] = 64'd0;
	mem_3[85] = 64'd0;
	mem_3[86] = 64'd0;
	mem_3[87] = 64'd0;
	mem_3[88] = 64'd0;
	mem_3[89] = 64'd0;
	mem_3[90] = 64'd0;
	mem_3[91] = 64'd0;
	mem_3[92] = 64'd0;
	mem_3[93] = 64'd0;
	mem_3[94] = 64'd0;
	mem_3[95] = 64'd0;
	mem_3[96] = 64'd0;
	mem_3[97] = 64'd0;
	mem_3[98] = 64'd0;
	mem_3[99] = 64'd0;
	mem_3[100] = 64'd0;
	mem_3[101] = 64'd0;
	mem_3[102] = 64'd0;
	mem_3[103] = 64'd0;
	mem_3[104] = 64'd0;
	mem_3[105] = 64'd0;
	mem_3[106] = 64'd0;
	mem_3[107] = 64'd0;
	mem_3[108] = 64'd0;
	mem_3[109] = 64'd0;
	mem_3[110] = 64'd0;
	mem_3[111] = 64'd0;
	mem_3[112] = 64'd0;
	mem_3[113] = 64'd0;
	mem_3[114] = 64'd0;
	mem_3[115] = 64'd0;
	mem_3[116] = 64'd0;
	mem_3[117] = 64'd0;
	mem_3[118] = 64'd0;
	mem_3[119] = 64'd0;
	mem_3[120] = 64'd0;
	mem_3[121] = 64'd0;
	mem_3[122] = 64'd0;
	mem_3[123] = 64'd0;
	mem_3[124] = 64'd0;
	mem_3[125] = 64'd0;
	mem_3[126] = 64'd0;
	mem_3[127] = 64'd0;
	mem_3[128] = 64'd0;
	mem_3[129] = 64'd0;
	mem_3[130] = 64'd0;
	mem_3[131] = 64'd0;
	mem_3[132] = 64'd0;
	mem_3[133] = 64'd0;
	mem_3[134] = 64'd0;
	mem_3[135] = 64'd0;
	mem_3[136] = 64'd0;
	mem_3[137] = 64'd0;
	mem_3[138] = 64'd0;
	mem_3[139] = 64'd0;
	mem_3[140] = 64'd0;
	mem_3[141] = 64'd0;
	mem_3[142] = 64'd0;
	mem_3[143] = 64'd0;
	mem_3[144] = 64'd0;
	mem_3[145] = 64'd0;
	mem_3[146] = 64'd0;
	mem_3[147] = 64'd0;
	mem_3[148] = 64'd0;
	mem_3[149] = 64'd0;
	mem_3[150] = 64'd0;
	mem_3[151] = 64'd0;
	mem_3[152] = 64'd0;
	mem_3[153] = 64'd0;
	mem_3[154] = 64'd0;
	mem_3[155] = 64'd0;
	mem_3[156] = 64'd0;
	mem_3[157] = 64'd0;
	mem_3[158] = 64'd0;
	mem_3[159] = 64'd0;
	mem_3[160] = 64'd0;
	mem_3[161] = 64'd0;
	mem_3[162] = 64'd0;
	mem_3[163] = 64'd0;
	mem_3[164] = 64'd0;
	mem_3[165] = 64'd0;
	mem_3[166] = 64'd0;
	mem_3[167] = 64'd0;
	mem_3[168] = 64'd0;
	mem_3[169] = 64'd0;
	mem_3[170] = 64'd0;
	mem_3[171] = 64'd0;
	mem_3[172] = 64'd0;
	mem_3[173] = 64'd0;
	mem_3[174] = 64'd0;
	mem_3[175] = 64'd0;
	mem_3[176] = 64'd0;
	mem_3[177] = 64'd0;
	mem_3[178] = 64'd0;
	mem_3[179] = 64'd0;
	mem_3[180] = 64'd0;
	mem_3[181] = 64'd0;
	mem_3[182] = 64'd0;
	mem_3[183] = 64'd0;
	mem_3[184] = 64'd0;
	mem_3[185] = 64'd0;
	mem_3[186] = 64'd0;
	mem_3[187] = 64'd0;
	mem_3[188] = 64'd0;
	mem_3[189] = 64'd0;
	mem_3[190] = 64'd0;
	mem_3[191] = 64'd0;
	mem_3[192] = 64'd0;
	mem_3[193] = 64'd0;
	mem_3[194] = 64'd0;
	mem_3[195] = 64'd0;
	mem_3[196] = 64'd0;
	mem_3[197] = 64'd0;
	mem_3[198] = 64'd0;
	mem_3[199] = 64'd0;
	mem_3[200] = 64'd0;
	mem_3[201] = 64'd0;
	mem_3[202] = 64'd0;
	mem_3[203] = 64'd0;
	mem_3[204] = 64'd0;
	mem_3[205] = 64'd0;
	mem_3[206] = 64'd0;
	mem_3[207] = 64'd0;
	mem_3[208] = 64'd0;
	mem_3[209] = 64'd0;
	mem_3[210] = 64'd0;
	mem_3[211] = 64'd0;
	mem_3[212] = 64'd0;
	mem_3[213] = 64'd0;
	mem_3[214] = 64'd0;
	mem_3[215] = 64'd0;
	mem_3[216] = 64'd0;
	mem_3[217] = 64'd0;
	mem_3[218] = 64'd0;
	mem_3[219] = 64'd0;
	mem_3[220] = 64'd0;
	mem_3[221] = 64'd0;
	mem_3[222] = 64'd0;
	mem_3[223] = 64'd0;
	mem_3[224] = 64'd0;
	mem_3[225] = 64'd0;
	mem_3[226] = 64'd0;
	mem_3[227] = 64'd0;
	mem_3[228] = 64'd0;
	mem_3[229] = 64'd0;
	mem_3[230] = 64'd0;
	mem_3[231] = 64'd0;
	mem_3[232] = 64'd0;
	mem_3[233] = 64'd0;
	mem_3[234] = 64'd0;
	mem_3[235] = 64'd0;
	mem_3[236] = 64'd0;
	mem_3[237] = 64'd0;
	mem_3[238] = 64'd0;
	mem_3[239] = 64'd0;
	mem_3[240] = 64'd0;
	mem_3[241] = 64'd0;
	mem_3[242] = 64'd0;
	mem_3[243] = 64'd0;
	mem_3[244] = 64'd0;
	mem_3[245] = 64'd0;
	mem_3[246] = 64'd0;
	mem_3[247] = 64'd0;
	mem_3[248] = 64'd0;
	mem_3[249] = 64'd0;
	mem_3[250] = 64'd0;
	mem_3[251] = 64'd0;
	mem_3[252] = 64'd0;
	mem_3[253] = 64'd0;
	mem_3[254] = 64'd0;
	mem_3[255] = 64'd0;
	mem_3[256] = 64'd0;
	mem_3[257] = 64'd0;
	mem_3[258] = 64'd0;
	mem_3[259] = 64'd0;
	mem_3[260] = 64'd0;
	mem_3[261] = 64'd0;
	mem_3[262] = 64'd0;
	mem_3[263] = 64'd0;
	mem_3[264] = 64'd0;
	mem_3[265] = 64'd0;
	mem_3[266] = 64'd0;
	mem_3[267] = 64'd0;
	mem_3[268] = 64'd0;
	mem_3[269] = 64'd0;
	mem_3[270] = 64'd0;
	mem_3[271] = 64'd0;
	mem_3[272] = 64'd0;
	mem_3[273] = 64'd0;
	mem_3[274] = 64'd0;
	mem_3[275] = 64'd0;
	mem_3[276] = 64'd0;
	mem_3[277] = 64'd0;
	mem_3[278] = 64'd0;
	mem_3[279] = 64'd0;
	mem_3[280] = 64'd0;
	mem_3[281] = 64'd0;
	mem_3[282] = 64'd0;
	mem_3[283] = 64'd0;
	mem_3[284] = 64'd0;
	mem_3[285] = 64'd0;
	mem_3[286] = 64'd0;
	mem_3[287] = 64'd0;
	mem_3[288] = 64'd0;
	mem_3[289] = 64'd0;
	mem_3[290] = 64'd0;
	mem_3[291] = 64'd0;
	mem_3[292] = 64'd0;
	mem_3[293] = 64'd0;
	mem_3[294] = 64'd0;
	mem_3[295] = 64'd0;
	mem_3[296] = 64'd0;
	mem_3[297] = 64'd0;
	mem_3[298] = 64'd0;
	mem_3[299] = 64'd0;
	mem_3[300] = 64'd0;
	mem_3[301] = 64'd0;
	mem_3[302] = 64'd0;
	mem_3[303] = 64'd0;
	mem_3[304] = 64'd0;
	mem_3[305] = 64'd0;
	mem_3[306] = 64'd0;
	mem_3[307] = 64'd0;
	mem_3[308] = 64'd0;
	mem_3[309] = 64'd0;
	mem_3[310] = 64'd0;
	mem_3[311] = 64'd0;
	mem_3[312] = 64'd0;
	mem_3[313] = 64'd0;
	mem_3[314] = 64'd0;
	mem_3[315] = 64'd0;
	mem_3[316] = 64'd0;
	mem_3[317] = 64'd0;
	mem_3[318] = 64'd0;
	mem_3[319] = 64'd0;
	mem_3[320] = 64'd0;
	mem_3[321] = 64'd0;
	mem_3[322] = 64'd0;
	mem_3[323] = 64'd0;
	mem_3[324] = 64'd0;
	mem_3[325] = 64'd0;
	mem_3[326] = 64'd0;
	mem_3[327] = 64'd0;
	mem_3[328] = 64'd0;
	mem_3[329] = 64'd0;
	mem_3[330] = 64'd0;
	mem_3[331] = 64'd0;
	mem_3[332] = 64'd0;
	mem_3[333] = 64'd0;
	mem_3[334] = 64'd0;
	mem_3[335] = 64'd0;
	mem_3[336] = 64'd0;
	mem_3[337] = 64'd0;
	mem_3[338] = 64'd0;
	mem_3[339] = 64'd0;
	mem_3[340] = 64'd0;
	mem_3[341] = 64'd0;
	mem_3[342] = 64'd0;
	mem_3[343] = 64'd0;
	mem_3[344] = 64'd0;
	mem_3[345] = 64'd0;
	mem_3[346] = 64'd0;
	mem_3[347] = 64'd0;
	mem_3[348] = 64'd0;
	mem_3[349] = 64'd0;
	mem_3[350] = 64'd0;
	mem_3[351] = 64'd0;
	mem_3[352] = 64'd0;
	mem_3[353] = 64'd0;
	mem_3[354] = 64'd0;
	mem_3[355] = 64'd0;
	mem_3[356] = 64'd0;
	mem_3[357] = 64'd0;
	mem_3[358] = 64'd0;
	mem_3[359] = 64'd0;
	mem_3[360] = 64'd0;
	mem_3[361] = 64'd0;
	mem_3[362] = 64'd0;
	mem_3[363] = 64'd0;
	mem_3[364] = 64'd0;
	mem_3[365] = 64'd0;
	mem_3[366] = 64'd0;
	mem_3[367] = 64'd0;
	mem_3[368] = 64'd0;
	mem_3[369] = 64'd0;
	mem_3[370] = 64'd0;
	mem_3[371] = 64'd0;
	mem_3[372] = 64'd0;
	mem_3[373] = 64'd0;
	mem_3[374] = 64'd0;
	mem_3[375] = 64'd0;
	mem_3[376] = 64'd0;
	mem_3[377] = 64'd0;
	mem_3[378] = 64'd0;
	mem_3[379] = 64'd0;
	mem_3[380] = 64'd0;
	mem_3[381] = 64'd0;
	mem_3[382] = 64'd0;
	mem_3[383] = 64'd0;
	mem_3[384] = 64'd0;
	mem_3[385] = 64'd0;
	mem_3[386] = 64'd0;
	mem_3[387] = 64'd0;
	mem_3[388] = 64'd0;
	mem_3[389] = 64'd0;
	mem_3[390] = 64'd0;
	mem_3[391] = 64'd0;
	mem_3[392] = 64'd0;
	mem_3[393] = 64'd0;
	mem_3[394] = 64'd0;
	mem_3[395] = 64'd0;
	mem_3[396] = 64'd0;
	mem_3[397] = 64'd0;
	mem_3[398] = 64'd0;
	mem_3[399] = 64'd0;
	mem_3[400] = 64'd0;
	mem_3[401] = 64'd0;
	mem_3[402] = 64'd0;
	mem_3[403] = 64'd0;
	mem_3[404] = 64'd0;
	mem_3[405] = 64'd0;
	mem_3[406] = 64'd0;
	mem_3[407] = 64'd0;
	mem_3[408] = 64'd0;
	mem_3[409] = 64'd0;
	mem_3[410] = 64'd0;
	mem_3[411] = 64'd0;
	mem_3[412] = 64'd0;
	mem_3[413] = 64'd0;
	mem_3[414] = 64'd0;
	mem_3[415] = 64'd0;
	mem_3[416] = 64'd0;
	mem_3[417] = 64'd0;
	mem_3[418] = 64'd0;
	mem_3[419] = 64'd0;
	mem_3[420] = 64'd0;
	mem_3[421] = 64'd0;
	mem_3[422] = 64'd0;
	mem_3[423] = 64'd0;
	mem_3[424] = 64'd0;
	mem_3[425] = 64'd0;
	mem_3[426] = 64'd0;
	mem_3[427] = 64'd0;
	mem_3[428] = 64'd0;
	mem_3[429] = 64'd0;
	mem_3[430] = 64'd0;
	mem_3[431] = 64'd0;
	mem_3[432] = 64'd0;
	mem_3[433] = 64'd0;
	mem_3[434] = 64'd0;
	mem_3[435] = 64'd0;
	mem_3[436] = 64'd0;
	mem_3[437] = 64'd0;
	mem_3[438] = 64'd0;
	mem_3[439] = 64'd0;
	mem_3[440] = 64'd0;
	mem_3[441] = 64'd0;
	mem_3[442] = 64'd0;
	mem_3[443] = 64'd0;
	mem_3[444] = 64'd0;
	mem_3[445] = 64'd0;
	mem_3[446] = 64'd0;
	mem_3[447] = 64'd0;
	mem_3[448] = 64'd0;
	mem_3[449] = 64'd0;
	mem_3[450] = 64'd0;
	mem_3[451] = 64'd0;
	mem_3[452] = 64'd0;
	mem_3[453] = 64'd0;
	mem_3[454] = 64'd0;
	mem_3[455] = 64'd0;
	mem_3[456] = 64'd0;
	mem_3[457] = 64'd0;
	mem_3[458] = 64'd0;
	mem_3[459] = 64'd0;
	mem_3[460] = 64'd0;
	mem_3[461] = 64'd0;
	mem_3[462] = 64'd0;
	mem_3[463] = 64'd0;
	mem_3[464] = 64'd0;
	mem_3[465] = 64'd0;
	mem_3[466] = 64'd0;
	mem_3[467] = 64'd0;
	mem_3[468] = 64'd0;
	mem_3[469] = 64'd0;
	mem_3[470] = 64'd0;
	mem_3[471] = 64'd0;
	mem_3[472] = 64'd0;
	mem_3[473] = 64'd0;
	mem_3[474] = 64'd0;
	mem_3[475] = 64'd0;
	mem_3[476] = 64'd0;
	mem_3[477] = 64'd0;
	mem_3[478] = 64'd0;
	mem_3[479] = 64'd0;
	mem_3[480] = 64'd0;
	mem_3[481] = 64'd0;
	mem_3[482] = 64'd0;
	mem_3[483] = 64'd0;
	mem_3[484] = 64'd0;
	mem_3[485] = 64'd0;
	mem_3[486] = 64'd0;
	mem_3[487] = 64'd0;
	mem_3[488] = 64'd0;
	mem_3[489] = 64'd0;
	mem_3[490] = 64'd0;
	mem_3[491] = 64'd0;
	mem_3[492] = 64'd0;
	mem_3[493] = 64'd0;
	mem_3[494] = 64'd0;
	mem_3[495] = 64'd0;
	mem_3[496] = 64'd0;
	mem_3[497] = 64'd0;
	mem_3[498] = 64'd0;
	mem_3[499] = 64'd0;
	mem_3[500] = 64'd0;
	mem_3[501] = 64'd0;
	mem_3[502] = 64'd0;
	mem_3[503] = 64'd0;
	mem_3[504] = 64'd0;
	mem_3[505] = 64'd0;
	mem_3[506] = 64'd0;
	mem_3[507] = 64'd0;
	mem_3[508] = 64'd0;
	mem_3[509] = 64'd0;
	mem_3[510] = 64'd0;
	mem_3[511] = 64'd0;
	mem_3[512] = 64'd0;
	mem_3[513] = 64'd0;
	mem_3[514] = 64'd0;
	mem_3[515] = 64'd0;
	mem_3[516] = 64'd0;
	mem_3[517] = 64'd0;
	mem_3[518] = 64'd0;
	mem_3[519] = 64'd0;
	mem_3[520] = 64'd0;
	mem_3[521] = 64'd0;
	mem_3[522] = 64'd0;
	mem_3[523] = 64'd0;
	mem_3[524] = 64'd0;
	mem_3[525] = 64'd0;
	mem_3[526] = 64'd0;
	mem_3[527] = 64'd0;
	mem_3[528] = 64'd0;
	mem_3[529] = 64'd0;
	mem_3[530] = 64'd0;
	mem_3[531] = 64'd0;
	mem_3[532] = 64'd0;
	mem_3[533] = 64'd0;
	mem_3[534] = 64'd0;
	mem_3[535] = 64'd0;
	mem_3[536] = 64'd0;
	mem_3[537] = 64'd0;
	mem_3[538] = 64'd0;
	mem_3[539] = 64'd0;
	mem_3[540] = 64'd0;
	mem_3[541] = 64'd0;
	mem_3[542] = 64'd0;
	mem_3[543] = 64'd0;
	mem_3[544] = 64'd0;
	mem_3[545] = 64'd0;
	mem_3[546] = 64'd0;
	mem_3[547] = 64'd0;
	mem_3[548] = 64'd0;
	mem_3[549] = 64'd0;
	mem_3[550] = 64'd0;
	mem_3[551] = 64'd0;
	mem_3[552] = 64'd0;
	mem_3[553] = 64'd0;
	mem_3[554] = 64'd0;
	mem_3[555] = 64'd0;
	mem_3[556] = 64'd0;
	mem_3[557] = 64'd0;
	mem_3[558] = 64'd0;
	mem_3[559] = 64'd0;
	mem_3[560] = 64'd0;
	mem_3[561] = 64'd0;
	mem_3[562] = 64'd0;
	mem_3[563] = 64'd0;
	mem_3[564] = 64'd0;
	mem_3[565] = 64'd0;
	mem_3[566] = 64'd0;
	mem_3[567] = 64'd0;
	mem_3[568] = 64'd0;
	mem_3[569] = 64'd0;
	mem_3[570] = 64'd0;
	mem_3[571] = 64'd0;
	mem_3[572] = 64'd0;
	mem_3[573] = 64'd0;
	mem_3[574] = 64'd0;
	mem_3[575] = 64'd0;
	mem_3[576] = 64'd0;
	mem_3[577] = 64'd0;
	mem_3[578] = 64'd0;
	mem_3[579] = 64'd0;
	mem_3[580] = 64'd0;
	mem_3[581] = 64'd0;
	mem_3[582] = 64'd0;
	mem_3[583] = 64'd0;
	mem_3[584] = 64'd0;
	mem_3[585] = 64'd0;
	mem_3[586] = 64'd0;
	mem_3[587] = 64'd0;
	mem_3[588] = 64'd0;
	mem_3[589] = 64'd0;
	mem_3[590] = 64'd0;
	mem_3[591] = 64'd0;
	mem_3[592] = 64'd0;
	mem_3[593] = 64'd0;
	mem_3[594] = 64'd0;
	mem_3[595] = 64'd0;
	mem_3[596] = 64'd0;
	mem_3[597] = 64'd0;
	mem_3[598] = 64'd0;
	mem_3[599] = 64'd0;
	mem_3[600] = 64'd0;
	mem_3[601] = 64'd0;
	mem_3[602] = 64'd0;
	mem_3[603] = 64'd0;
	mem_3[604] = 64'd0;
	mem_3[605] = 64'd0;
	mem_3[606] = 64'd0;
	mem_3[607] = 64'd0;
	mem_3[608] = 64'd0;
	mem_3[609] = 64'd0;
	mem_3[610] = 64'd0;
	mem_3[611] = 64'd0;
	mem_3[612] = 64'd0;
	mem_3[613] = 64'd0;
	mem_3[614] = 64'd0;
	mem_3[615] = 64'd0;
	mem_3[616] = 64'd0;
	mem_3[617] = 64'd0;
	mem_3[618] = 64'd0;
	mem_3[619] = 64'd0;
	mem_3[620] = 64'd0;
	mem_3[621] = 64'd0;
	mem_3[622] = 64'd0;
	mem_3[623] = 64'd0;
	mem_3[624] = 64'd0;
	mem_3[625] = 64'd0;
	mem_3[626] = 64'd0;
	mem_3[627] = 64'd0;
	mem_3[628] = 64'd0;
	mem_3[629] = 64'd0;
	mem_3[630] = 64'd0;
	mem_3[631] = 64'd0;
	mem_3[632] = 64'd0;
	mem_3[633] = 64'd0;
	mem_3[634] = 64'd0;
	mem_3[635] = 64'd0;
	mem_3[636] = 64'd0;
	mem_3[637] = 64'd0;
	mem_3[638] = 64'd0;
	mem_3[639] = 64'd0;
	mem_3[640] = 64'd0;
	mem_3[641] = 64'd0;
	mem_3[642] = 64'd0;
	mem_3[643] = 64'd0;
	mem_3[644] = 64'd0;
	mem_3[645] = 64'd0;
	mem_3[646] = 64'd0;
	mem_3[647] = 64'd0;
	mem_3[648] = 64'd0;
	mem_3[649] = 64'd0;
	mem_3[650] = 64'd0;
	mem_3[651] = 64'd0;
	mem_3[652] = 64'd0;
	mem_3[653] = 64'd0;
	mem_3[654] = 64'd0;
	mem_3[655] = 64'd0;
	mem_3[656] = 64'd0;
	mem_3[657] = 64'd0;
	mem_3[658] = 64'd0;
	mem_3[659] = 64'd0;
	mem_3[660] = 64'd0;
	mem_3[661] = 64'd0;
	mem_3[662] = 64'd0;
	mem_3[663] = 64'd0;
	mem_3[664] = 64'd0;
	mem_3[665] = 64'd0;
	mem_3[666] = 64'd0;
	mem_3[667] = 64'd0;
	mem_3[668] = 64'd0;
	mem_3[669] = 64'd0;
	mem_3[670] = 64'd0;
	mem_3[671] = 64'd0;
	mem_3[672] = 64'd0;
	mem_3[673] = 64'd0;
	mem_3[674] = 64'd0;
	mem_3[675] = 64'd0;
	mem_3[676] = 64'd0;
	mem_3[677] = 64'd0;
	mem_3[678] = 64'd0;
	mem_3[679] = 64'd0;
	mem_3[680] = 64'd0;
	mem_3[681] = 64'd0;
	mem_3[682] = 64'd0;
	mem_3[683] = 64'd0;
	mem_3[684] = 64'd0;
	mem_3[685] = 64'd0;
	mem_3[686] = 64'd0;
	mem_3[687] = 64'd0;
	mem_3[688] = 64'd0;
	mem_3[689] = 64'd0;
	mem_3[690] = 64'd0;
	mem_3[691] = 64'd0;
	mem_3[692] = 64'd0;
	mem_3[693] = 64'd0;
	mem_3[694] = 64'd0;
	mem_3[695] = 64'd0;
	mem_3[696] = 64'd0;
	mem_3[697] = 64'd0;
	mem_3[698] = 64'd0;
	mem_3[699] = 64'd0;
	mem_3[700] = 64'd0;
	mem_3[701] = 64'd0;
	mem_3[702] = 64'd0;
	mem_3[703] = 64'd0;
	mem_3[704] = 64'd0;
	mem_3[705] = 64'd0;
	mem_3[706] = 64'd0;
	mem_3[707] = 64'd0;
	mem_3[708] = 64'd0;
	mem_3[709] = 64'd0;
	mem_3[710] = 64'd0;
	mem_3[711] = 64'd0;
	mem_3[712] = 64'd0;
	mem_3[713] = 64'd0;
	mem_3[714] = 64'd0;
	mem_3[715] = 64'd0;
	mem_3[716] = 64'd0;
	mem_3[717] = 64'd0;
	mem_3[718] = 64'd0;
	mem_3[719] = 64'd0;
	mem_3[720] = 64'd0;
	mem_3[721] = 64'd0;
	mem_3[722] = 64'd0;
	mem_3[723] = 64'd0;
	mem_3[724] = 64'd0;
	mem_3[725] = 64'd0;
	mem_3[726] = 64'd0;
	mem_3[727] = 64'd0;
	mem_3[728] = 64'd0;
	mem_3[729] = 64'd0;
	mem_3[730] = 64'd0;
	mem_3[731] = 64'd0;
	mem_3[732] = 64'd0;
	mem_3[733] = 64'd0;
	mem_3[734] = 64'd0;
	mem_3[735] = 64'd0;
	mem_3[736] = 64'd0;
	mem_3[737] = 64'd0;
	mem_3[738] = 64'd0;
	mem_3[739] = 64'd0;
	mem_3[740] = 64'd0;
	mem_3[741] = 64'd0;
	mem_3[742] = 64'd0;
	mem_3[743] = 64'd0;
	mem_3[744] = 64'd0;
	mem_3[745] = 64'd0;
	mem_3[746] = 64'd0;
	mem_3[747] = 64'd0;
	mem_3[748] = 64'd0;
	mem_3[749] = 64'd0;
	mem_3[750] = 64'd0;
	mem_3[751] = 64'd0;
	mem_3[752] = 64'd0;
	mem_3[753] = 64'd0;
	mem_3[754] = 64'd0;
	mem_3[755] = 64'd0;
	mem_3[756] = 64'd0;
	mem_3[757] = 64'd0;
	mem_3[758] = 64'd0;
	mem_3[759] = 64'd0;
	mem_3[760] = 64'd0;
	mem_3[761] = 64'd0;
	mem_3[762] = 64'd0;
	mem_3[763] = 64'd0;
	mem_3[764] = 64'd0;
	mem_3[765] = 64'd0;
	mem_3[766] = 64'd0;
	mem_3[767] = 64'd0;
	mem_3[768] = 64'd0;
	mem_3[769] = 64'd0;
	mem_3[770] = 64'd0;
	mem_3[771] = 64'd0;
	mem_3[772] = 64'd0;
	mem_3[773] = 64'd0;
	mem_3[774] = 64'd0;
	mem_3[775] = 64'd0;
	mem_3[776] = 64'd0;
	mem_3[777] = 64'd0;
	mem_3[778] = 64'd0;
	mem_3[779] = 64'd0;
	mem_3[780] = 64'd0;
	mem_3[781] = 64'd0;
	mem_3[782] = 64'd0;
	mem_3[783] = 64'd0;
	mem_3[784] = 64'd0;
	mem_3[785] = 64'd0;
	mem_3[786] = 64'd0;
	mem_3[787] = 64'd0;
	mem_3[788] = 64'd0;
	mem_3[789] = 64'd0;
	mem_3[790] = 64'd0;
	mem_3[791] = 64'd0;
	mem_3[792] = 64'd0;
	mem_3[793] = 64'd0;
	mem_3[794] = 64'd0;
	mem_3[795] = 64'd0;
	mem_3[796] = 64'd0;
	mem_3[797] = 64'd0;
	mem_3[798] = 64'd0;
	mem_3[799] = 64'd0;
	mem_3[800] = 64'd0;
	mem_3[801] = 64'd0;
	mem_3[802] = 64'd0;
	mem_3[803] = 64'd0;
	mem_3[804] = 64'd0;
	mem_3[805] = 64'd0;
	mem_3[806] = 64'd0;
	mem_3[807] = 64'd0;
	mem_3[808] = 64'd0;
	mem_3[809] = 64'd0;
	mem_3[810] = 64'd0;
	mem_3[811] = 64'd0;
	mem_3[812] = 64'd0;
	mem_3[813] = 64'd0;
	mem_3[814] = 64'd0;
	mem_3[815] = 64'd0;
	mem_3[816] = 64'd0;
	mem_3[817] = 64'd0;
	mem_3[818] = 64'd0;
	mem_3[819] = 64'd0;
	mem_3[820] = 64'd0;
	mem_3[821] = 64'd0;
	mem_3[822] = 64'd0;
	mem_3[823] = 64'd0;
	mem_3[824] = 64'd0;
	mem_3[825] = 64'd0;
	mem_3[826] = 64'd0;
	mem_3[827] = 64'd0;
	mem_3[828] = 64'd0;
	mem_3[829] = 64'd0;
	mem_3[830] = 64'd0;
	mem_3[831] = 64'd0;
	mem_3[832] = 64'd0;
	mem_3[833] = 64'd0;
	mem_3[834] = 64'd0;
	mem_3[835] = 64'd0;
	mem_3[836] = 64'd0;
	mem_3[837] = 64'd0;
	mem_3[838] = 64'd0;
	mem_3[839] = 64'd0;
	mem_3[840] = 64'd0;
	mem_3[841] = 64'd0;
	mem_3[842] = 64'd0;
	mem_3[843] = 64'd0;
	mem_3[844] = 64'd0;
	mem_3[845] = 64'd0;
	mem_3[846] = 64'd0;
	mem_3[847] = 64'd0;
	mem_3[848] = 64'd0;
	mem_3[849] = 64'd0;
	mem_3[850] = 64'd0;
	mem_3[851] = 64'd0;
	mem_3[852] = 64'd0;
	mem_3[853] = 64'd0;
	mem_3[854] = 64'd0;
	mem_3[855] = 64'd0;
	mem_3[856] = 64'd0;
	mem_3[857] = 64'd0;
	mem_3[858] = 64'd0;
	mem_3[859] = 64'd0;
	mem_3[860] = 64'd0;
	mem_3[861] = 64'd0;
	mem_3[862] = 64'd0;
	mem_3[863] = 64'd0;
	mem_3[864] = 64'd0;
	mem_3[865] = 64'd0;
	mem_3[866] = 64'd0;
	mem_3[867] = 64'd0;
	mem_3[868] = 64'd0;
	mem_3[869] = 64'd0;
	mem_3[870] = 64'd0;
	mem_3[871] = 64'd0;
	mem_3[872] = 64'd0;
	mem_3[873] = 64'd0;
	mem_3[874] = 64'd0;
	mem_3[875] = 64'd0;
	mem_3[876] = 64'd0;
	mem_3[877] = 64'd0;
	mem_3[878] = 64'd0;
	mem_3[879] = 64'd0;
	mem_3[880] = 64'd0;
	mem_3[881] = 64'd0;
	mem_3[882] = 64'd0;
	mem_3[883] = 64'd0;
	mem_3[884] = 64'd0;
	mem_3[885] = 64'd0;
	mem_3[886] = 64'd0;
	mem_3[887] = 64'd0;
	mem_3[888] = 64'd0;
	mem_3[889] = 64'd0;
	mem_3[890] = 64'd0;
	mem_3[891] = 64'd0;
	mem_3[892] = 64'd0;
	mem_3[893] = 64'd0;
	mem_3[894] = 64'd0;
	mem_3[895] = 64'd0;
	mem_3[896] = 64'd0;
	mem_3[897] = 64'd0;
	mem_3[898] = 64'd0;
	mem_3[899] = 64'd0;
	mem_3[900] = 64'd0;
	mem_3[901] = 64'd0;
	mem_3[902] = 64'd0;
	mem_3[903] = 64'd0;
	mem_3[904] = 64'd0;
	mem_3[905] = 64'd0;
	mem_3[906] = 64'd0;
	mem_3[907] = 64'd0;
	mem_3[908] = 64'd0;
	mem_3[909] = 64'd0;
	mem_3[910] = 64'd0;
	mem_3[911] = 64'd0;
	mem_3[912] = 64'd0;
	mem_3[913] = 64'd0;
	mem_3[914] = 64'd0;
	mem_3[915] = 64'd0;
	mem_3[916] = 64'd0;
	mem_3[917] = 64'd0;
	mem_3[918] = 64'd0;
	mem_3[919] = 64'd0;
	mem_3[920] = 64'd0;
	mem_3[921] = 64'd0;
	mem_3[922] = 64'd0;
	mem_3[923] = 64'd0;
	mem_3[924] = 64'd0;
	mem_3[925] = 64'd0;
	mem_3[926] = 64'd0;
	mem_3[927] = 64'd0;
	mem_3[928] = 64'd0;
	mem_3[929] = 64'd0;
	mem_3[930] = 64'd0;
	mem_3[931] = 64'd0;
	mem_3[932] = 64'd0;
	mem_3[933] = 64'd0;
	mem_3[934] = 64'd0;
	mem_3[935] = 64'd0;
	mem_3[936] = 64'd0;
	mem_3[937] = 64'd0;
	mem_3[938] = 64'd0;
	mem_3[939] = 64'd0;
	mem_3[940] = 64'd0;
	mem_3[941] = 64'd0;
	mem_3[942] = 64'd0;
	mem_3[943] = 64'd0;
	mem_3[944] = 64'd0;
	mem_3[945] = 64'd0;
	mem_3[946] = 64'd0;
	mem_3[947] = 64'd0;
	mem_3[948] = 64'd0;
	mem_3[949] = 64'd0;
	mem_3[950] = 64'd0;
	mem_3[951] = 64'd0;
	mem_3[952] = 64'd0;
	mem_3[953] = 64'd0;
	mem_3[954] = 64'd0;
	mem_3[955] = 64'd0;
	mem_3[956] = 64'd0;
	mem_3[957] = 64'd0;
	mem_3[958] = 64'd0;
	mem_3[959] = 64'd0;
	mem_3[960] = 64'd0;
	mem_3[961] = 64'd0;
	mem_3[962] = 64'd0;
	mem_3[963] = 64'd0;
	mem_3[964] = 64'd0;
	mem_3[965] = 64'd0;
	mem_3[966] = 64'd0;
	mem_3[967] = 64'd0;
	mem_3[968] = 64'd0;
	mem_3[969] = 64'd0;
	mem_3[970] = 64'd0;
	mem_3[971] = 64'd0;
	mem_3[972] = 64'd0;
	mem_3[973] = 64'd0;
	mem_3[974] = 64'd0;
	mem_3[975] = 64'd0;
	mem_3[976] = 64'd0;
	mem_3[977] = 64'd0;
	mem_3[978] = 64'd0;
	mem_3[979] = 64'd0;
	mem_3[980] = 64'd0;
	mem_3[981] = 64'd0;
	mem_3[982] = 64'd0;
	mem_3[983] = 64'd0;
	mem_3[984] = 64'd0;
	mem_3[985] = 64'd0;
	mem_3[986] = 64'd0;
	mem_3[987] = 64'd0;
	mem_3[988] = 64'd0;
	mem_3[989] = 64'd0;
	mem_3[990] = 64'd0;
	mem_3[991] = 64'd0;
	mem_3[992] = 64'd0;
	mem_3[993] = 64'd0;
	mem_3[994] = 64'd0;
	mem_3[995] = 64'd0;
	mem_3[996] = 64'd0;
	mem_3[997] = 64'd0;
	mem_3[998] = 64'd0;
	mem_3[999] = 64'd0;
	mem_3[1000] = 64'd0;
	mem_3[1001] = 64'd0;
	mem_3[1002] = 64'd0;
	mem_3[1003] = 64'd0;
	mem_3[1004] = 64'd0;
	mem_3[1005] = 64'd0;
	mem_3[1006] = 64'd0;
	mem_3[1007] = 64'd0;
	mem_3[1008] = 64'd0;
	mem_3[1009] = 64'd0;
	mem_3[1010] = 64'd0;
	mem_3[1011] = 64'd0;
	mem_3[1012] = 64'd0;
	mem_3[1013] = 64'd0;
	mem_3[1014] = 64'd0;
	mem_3[1015] = 64'd0;
	mem_3[1016] = 64'd0;
	mem_3[1017] = 64'd0;
	mem_3[1018] = 64'd0;
	mem_3[1019] = 64'd0;
	mem_3[1020] = 64'd0;
	mem_3[1021] = 64'd0;
	mem_3[1022] = 64'd0;
	mem_3[1023] = 64'd0;
	mem_4[0] = 64'd0;
	mem_4[1] = 64'd0;
	mem_4[2] = 64'd0;
	mem_4[3] = 64'd0;
	mem_4[4] = 64'd0;
	mem_4[5] = 64'd0;
	mem_4[6] = 64'd0;
	mem_4[7] = 64'd0;
	mem_4[8] = 64'd0;
	mem_4[9] = 64'd0;
	mem_4[10] = 64'd0;
	mem_4[11] = 64'd0;
	mem_4[12] = 64'd0;
	mem_4[13] = 64'd0;
	mem_4[14] = 64'd0;
	mem_4[15] = 64'd0;
	mem_4[16] = 64'd0;
	mem_4[17] = 64'd0;
	mem_4[18] = 64'd0;
	mem_4[19] = 64'd0;
	mem_4[20] = 64'd0;
	mem_4[21] = 64'd0;
	mem_4[22] = 64'd0;
	mem_4[23] = 64'd0;
	mem_4[24] = 64'd0;
	mem_4[25] = 64'd0;
	mem_4[26] = 64'd0;
	mem_4[27] = 64'd0;
	mem_4[28] = 64'd0;
	mem_4[29] = 64'd0;
	mem_4[30] = 64'd0;
	mem_4[31] = 64'd0;
	mem_4[32] = 64'd0;
	mem_4[33] = 64'd0;
	mem_4[34] = 64'd0;
	mem_4[35] = 64'd0;
	mem_4[36] = 64'd0;
	mem_4[37] = 64'd0;
	mem_4[38] = 64'd0;
	mem_4[39] = 64'd0;
	mem_4[40] = 64'd0;
	mem_4[41] = 64'd0;
	mem_4[42] = 64'd0;
	mem_4[43] = 64'd0;
	mem_4[44] = 64'd0;
	mem_4[45] = 64'd0;
	mem_4[46] = 64'd0;
	mem_4[47] = 64'd0;
	mem_4[48] = 64'd0;
	mem_4[49] = 64'd0;
	mem_4[50] = 64'd0;
	mem_4[51] = 64'd0;
	mem_4[52] = 64'd0;
	mem_4[53] = 64'd0;
	mem_4[54] = 64'd0;
	mem_4[55] = 64'd0;
	mem_4[56] = 64'd0;
	mem_4[57] = 64'd0;
	mem_4[58] = 64'd0;
	mem_4[59] = 64'd0;
	mem_4[60] = 64'd0;
	mem_4[61] = 64'd0;
	mem_4[62] = 64'd0;
	mem_4[63] = 64'd0;
	mem_4[64] = 64'd0;
	mem_4[65] = 64'd0;
	mem_4[66] = 64'd0;
	mem_4[67] = 64'd0;
	mem_4[68] = 64'd0;
	mem_4[69] = 64'd0;
	mem_4[70] = 64'd0;
	mem_4[71] = 64'd0;
	mem_4[72] = 64'd0;
	mem_4[73] = 64'd0;
	mem_4[74] = 64'd0;
	mem_4[75] = 64'd0;
	mem_4[76] = 64'd0;
	mem_4[77] = 64'd0;
	mem_4[78] = 64'd0;
	mem_4[79] = 64'd0;
	mem_4[80] = 64'd0;
	mem_4[81] = 64'd0;
	mem_4[82] = 64'd0;
	mem_4[83] = 64'd0;
	mem_4[84] = 64'd0;
	mem_4[85] = 64'd0;
	mem_4[86] = 64'd0;
	mem_4[87] = 64'd0;
	mem_4[88] = 64'd0;
	mem_4[89] = 64'd0;
	mem_4[90] = 64'd0;
	mem_4[91] = 64'd0;
	mem_4[92] = 64'd0;
	mem_4[93] = 64'd0;
	mem_4[94] = 64'd0;
	mem_4[95] = 64'd0;
	mem_4[96] = 64'd0;
	mem_4[97] = 64'd0;
	mem_4[98] = 64'd0;
	mem_4[99] = 64'd0;
	mem_4[100] = 64'd0;
	mem_4[101] = 64'd0;
	mem_4[102] = 64'd0;
	mem_4[103] = 64'd0;
	mem_4[104] = 64'd0;
	mem_4[105] = 64'd0;
	mem_4[106] = 64'd0;
	mem_4[107] = 64'd0;
	mem_4[108] = 64'd0;
	mem_4[109] = 64'd0;
	mem_4[110] = 64'd0;
	mem_4[111] = 64'd0;
	mem_4[112] = 64'd0;
	mem_4[113] = 64'd0;
	mem_4[114] = 64'd0;
	mem_4[115] = 64'd0;
	mem_4[116] = 64'd0;
	mem_4[117] = 64'd0;
	mem_4[118] = 64'd0;
	mem_4[119] = 64'd0;
	mem_4[120] = 64'd0;
	mem_4[121] = 64'd0;
	mem_4[122] = 64'd0;
	mem_4[123] = 64'd0;
	mem_4[124] = 64'd0;
	mem_4[125] = 64'd0;
	mem_4[126] = 64'd0;
	mem_4[127] = 64'd0;
	mem_4[128] = 64'd0;
	mem_4[129] = 64'd0;
	mem_4[130] = 64'd0;
	mem_4[131] = 64'd0;
	mem_4[132] = 64'd0;
	mem_4[133] = 64'd0;
	mem_4[134] = 64'd0;
	mem_4[135] = 64'd0;
	mem_4[136] = 64'd0;
	mem_4[137] = 64'd0;
	mem_4[138] = 64'd0;
	mem_4[139] = 64'd0;
	mem_4[140] = 64'd0;
	mem_4[141] = 64'd0;
	mem_4[142] = 64'd0;
	mem_4[143] = 64'd0;
	mem_4[144] = 64'd0;
	mem_4[145] = 64'd0;
	mem_4[146] = 64'd0;
	mem_4[147] = 64'd0;
	mem_4[148] = 64'd0;
	mem_4[149] = 64'd0;
	mem_4[150] = 64'd0;
	mem_4[151] = 64'd0;
	mem_4[152] = 64'd0;
	mem_4[153] = 64'd0;
	mem_4[154] = 64'd0;
	mem_4[155] = 64'd0;
	mem_4[156] = 64'd0;
	mem_4[157] = 64'd0;
	mem_4[158] = 64'd0;
	mem_4[159] = 64'd0;
	mem_4[160] = 64'd0;
	mem_4[161] = 64'd0;
	mem_4[162] = 64'd0;
	mem_4[163] = 64'd0;
	mem_4[164] = 64'd0;
	mem_4[165] = 64'd0;
	mem_4[166] = 64'd0;
	mem_4[167] = 64'd0;
	mem_4[168] = 64'd0;
	mem_4[169] = 64'd0;
	mem_4[170] = 64'd0;
	mem_4[171] = 64'd0;
	mem_4[172] = 64'd0;
	mem_4[173] = 64'd0;
	mem_4[174] = 64'd0;
	mem_4[175] = 64'd0;
	mem_4[176] = 64'd0;
	mem_4[177] = 64'd0;
	mem_4[178] = 64'd0;
	mem_4[179] = 64'd0;
	mem_4[180] = 64'd0;
	mem_4[181] = 64'd0;
	mem_4[182] = 64'd0;
	mem_4[183] = 64'd0;
	mem_4[184] = 64'd0;
	mem_4[185] = 64'd0;
	mem_4[186] = 64'd0;
	mem_4[187] = 64'd0;
	mem_4[188] = 64'd0;
	mem_4[189] = 64'd0;
	mem_4[190] = 64'd0;
	mem_4[191] = 64'd0;
	mem_4[192] = 64'd0;
	mem_4[193] = 64'd0;
	mem_4[194] = 64'd0;
	mem_4[195] = 64'd0;
	mem_4[196] = 64'd0;
	mem_4[197] = 64'd0;
	mem_4[198] = 64'd0;
	mem_4[199] = 64'd0;
	mem_4[200] = 64'd0;
	mem_4[201] = 64'd0;
	mem_4[202] = 64'd0;
	mem_4[203] = 64'd0;
	mem_4[204] = 64'd0;
	mem_4[205] = 64'd0;
	mem_4[206] = 64'd0;
	mem_4[207] = 64'd0;
	mem_4[208] = 64'd0;
	mem_4[209] = 64'd0;
	mem_4[210] = 64'd0;
	mem_4[211] = 64'd0;
	mem_4[212] = 64'd0;
	mem_4[213] = 64'd0;
	mem_4[214] = 64'd0;
	mem_4[215] = 64'd0;
	mem_4[216] = 64'd0;
	mem_4[217] = 64'd0;
	mem_4[218] = 64'd0;
	mem_4[219] = 64'd0;
	mem_4[220] = 64'd0;
	mem_4[221] = 64'd0;
	mem_4[222] = 64'd0;
	mem_4[223] = 64'd0;
	mem_4[224] = 64'd0;
	mem_4[225] = 64'd0;
	mem_4[226] = 64'd0;
	mem_4[227] = 64'd0;
	mem_4[228] = 64'd0;
	mem_4[229] = 64'd0;
	mem_4[230] = 64'd0;
	mem_4[231] = 64'd0;
	mem_4[232] = 64'd0;
	mem_4[233] = 64'd0;
	mem_4[234] = 64'd0;
	mem_4[235] = 64'd0;
	mem_4[236] = 64'd0;
	mem_4[237] = 64'd0;
	mem_4[238] = 64'd0;
	mem_4[239] = 64'd0;
	mem_4[240] = 64'd0;
	mem_4[241] = 64'd0;
	mem_4[242] = 64'd0;
	mem_4[243] = 64'd0;
	mem_4[244] = 64'd0;
	mem_4[245] = 64'd0;
	mem_4[246] = 64'd0;
	mem_4[247] = 64'd0;
	mem_4[248] = 64'd0;
	mem_4[249] = 64'd0;
	mem_4[250] = 64'd0;
	mem_4[251] = 64'd0;
	mem_4[252] = 64'd0;
	mem_4[253] = 64'd0;
	mem_4[254] = 64'd0;
	mem_4[255] = 64'd0;
	mem_4[256] = 64'd0;
	mem_4[257] = 64'd0;
	mem_4[258] = 64'd0;
	mem_4[259] = 64'd0;
	mem_4[260] = 64'd0;
	mem_4[261] = 64'd0;
	mem_4[262] = 64'd0;
	mem_4[263] = 64'd0;
	mem_4[264] = 64'd0;
	mem_4[265] = 64'd0;
	mem_4[266] = 64'd0;
	mem_4[267] = 64'd0;
	mem_4[268] = 64'd0;
	mem_4[269] = 64'd0;
	mem_4[270] = 64'd0;
	mem_4[271] = 64'd0;
	mem_4[272] = 64'd0;
	mem_4[273] = 64'd0;
	mem_4[274] = 64'd0;
	mem_4[275] = 64'd0;
	mem_4[276] = 64'd0;
	mem_4[277] = 64'd0;
	mem_4[278] = 64'd0;
	mem_4[279] = 64'd0;
	mem_4[280] = 64'd0;
	mem_4[281] = 64'd0;
	mem_4[282] = 64'd0;
	mem_4[283] = 64'd0;
	mem_4[284] = 64'd0;
	mem_4[285] = 64'd0;
	mem_4[286] = 64'd0;
	mem_4[287] = 64'd0;
	mem_4[288] = 64'd0;
	mem_4[289] = 64'd0;
	mem_4[290] = 64'd0;
	mem_4[291] = 64'd0;
	mem_4[292] = 64'd0;
	mem_4[293] = 64'd0;
	mem_4[294] = 64'd0;
	mem_4[295] = 64'd0;
	mem_4[296] = 64'd0;
	mem_4[297] = 64'd0;
	mem_4[298] = 64'd0;
	mem_4[299] = 64'd0;
	mem_4[300] = 64'd0;
	mem_4[301] = 64'd0;
	mem_4[302] = 64'd0;
	mem_4[303] = 64'd0;
	mem_4[304] = 64'd0;
	mem_4[305] = 64'd0;
	mem_4[306] = 64'd0;
	mem_4[307] = 64'd0;
	mem_4[308] = 64'd0;
	mem_4[309] = 64'd0;
	mem_4[310] = 64'd0;
	mem_4[311] = 64'd0;
	mem_4[312] = 64'd0;
	mem_4[313] = 64'd0;
	mem_4[314] = 64'd0;
	mem_4[315] = 64'd0;
	mem_4[316] = 64'd0;
	mem_4[317] = 64'd0;
	mem_4[318] = 64'd0;
	mem_4[319] = 64'd0;
	mem_4[320] = 64'd0;
	mem_4[321] = 64'd0;
	mem_4[322] = 64'd0;
	mem_4[323] = 64'd0;
	mem_4[324] = 64'd0;
	mem_4[325] = 64'd0;
	mem_4[326] = 64'd0;
	mem_4[327] = 64'd0;
	mem_4[328] = 64'd0;
	mem_4[329] = 64'd0;
	mem_4[330] = 64'd0;
	mem_4[331] = 64'd0;
	mem_4[332] = 64'd0;
	mem_4[333] = 64'd0;
	mem_4[334] = 64'd0;
	mem_4[335] = 64'd0;
	mem_4[336] = 64'd0;
	mem_4[337] = 64'd0;
	mem_4[338] = 64'd0;
	mem_4[339] = 64'd0;
	mem_4[340] = 64'd0;
	mem_4[341] = 64'd0;
	mem_4[342] = 64'd0;
	mem_4[343] = 64'd0;
	mem_4[344] = 64'd0;
	mem_4[345] = 64'd0;
	mem_4[346] = 64'd0;
	mem_4[347] = 64'd0;
	mem_4[348] = 64'd0;
	mem_4[349] = 64'd0;
	mem_4[350] = 64'd0;
	mem_4[351] = 64'd0;
	mem_4[352] = 64'd0;
	mem_4[353] = 64'd0;
	mem_4[354] = 64'd0;
	mem_4[355] = 64'd0;
	mem_4[356] = 64'd0;
	mem_4[357] = 64'd0;
	mem_4[358] = 64'd0;
	mem_4[359] = 64'd0;
	mem_4[360] = 64'd0;
	mem_4[361] = 64'd0;
	mem_4[362] = 64'd0;
	mem_4[363] = 64'd0;
	mem_4[364] = 64'd0;
	mem_4[365] = 64'd0;
	mem_4[366] = 64'd0;
	mem_4[367] = 64'd0;
	mem_4[368] = 64'd0;
	mem_4[369] = 64'd0;
	mem_4[370] = 64'd0;
	mem_4[371] = 64'd0;
	mem_4[372] = 64'd0;
	mem_4[373] = 64'd0;
	mem_4[374] = 64'd0;
	mem_4[375] = 64'd0;
	mem_4[376] = 64'd0;
	mem_4[377] = 64'd0;
	mem_4[378] = 64'd0;
	mem_4[379] = 64'd0;
	mem_4[380] = 64'd0;
	mem_4[381] = 64'd0;
	mem_4[382] = 64'd0;
	mem_4[383] = 64'd0;
	mem_4[384] = 64'd0;
	mem_4[385] = 64'd0;
	mem_4[386] = 64'd0;
	mem_4[387] = 64'd0;
	mem_4[388] = 64'd0;
	mem_4[389] = 64'd0;
	mem_4[390] = 64'd0;
	mem_4[391] = 64'd0;
	mem_4[392] = 64'd0;
	mem_4[393] = 64'd0;
	mem_4[394] = 64'd0;
	mem_4[395] = 64'd0;
	mem_4[396] = 64'd0;
	mem_4[397] = 64'd0;
	mem_4[398] = 64'd0;
	mem_4[399] = 64'd0;
	mem_4[400] = 64'd0;
	mem_4[401] = 64'd0;
	mem_4[402] = 64'd0;
	mem_4[403] = 64'd0;
	mem_4[404] = 64'd0;
	mem_4[405] = 64'd0;
	mem_4[406] = 64'd0;
	mem_4[407] = 64'd0;
	mem_4[408] = 64'd0;
	mem_4[409] = 64'd0;
	mem_4[410] = 64'd0;
	mem_4[411] = 64'd0;
	mem_4[412] = 64'd0;
	mem_4[413] = 64'd0;
	mem_4[414] = 64'd0;
	mem_4[415] = 64'd0;
	mem_4[416] = 64'd0;
	mem_4[417] = 64'd0;
	mem_4[418] = 64'd0;
	mem_4[419] = 64'd0;
	mem_4[420] = 64'd0;
	mem_4[421] = 64'd0;
	mem_4[422] = 64'd0;
	mem_4[423] = 64'd0;
	mem_4[424] = 64'd0;
	mem_4[425] = 64'd0;
	mem_4[426] = 64'd0;
	mem_4[427] = 64'd0;
	mem_4[428] = 64'd0;
	mem_4[429] = 64'd0;
	mem_4[430] = 64'd0;
	mem_4[431] = 64'd0;
	mem_4[432] = 64'd0;
	mem_4[433] = 64'd0;
	mem_4[434] = 64'd0;
	mem_4[435] = 64'd0;
	mem_4[436] = 64'd0;
	mem_4[437] = 64'd0;
	mem_4[438] = 64'd0;
	mem_4[439] = 64'd0;
	mem_4[440] = 64'd0;
	mem_4[441] = 64'd0;
	mem_4[442] = 64'd0;
	mem_4[443] = 64'd0;
	mem_4[444] = 64'd0;
	mem_4[445] = 64'd0;
	mem_4[446] = 64'd0;
	mem_4[447] = 64'd0;
	mem_4[448] = 64'd0;
	mem_4[449] = 64'd0;
	mem_4[450] = 64'd0;
	mem_4[451] = 64'd0;
	mem_4[452] = 64'd0;
	mem_4[453] = 64'd0;
	mem_4[454] = 64'd0;
	mem_4[455] = 64'd0;
	mem_4[456] = 64'd0;
	mem_4[457] = 64'd0;
	mem_4[458] = 64'd0;
	mem_4[459] = 64'd0;
	mem_4[460] = 64'd0;
	mem_4[461] = 64'd0;
	mem_4[462] = 64'd0;
	mem_4[463] = 64'd0;
	mem_4[464] = 64'd0;
	mem_4[465] = 64'd0;
	mem_4[466] = 64'd0;
	mem_4[467] = 64'd0;
	mem_4[468] = 64'd0;
	mem_4[469] = 64'd0;
	mem_4[470] = 64'd0;
	mem_4[471] = 64'd0;
	mem_4[472] = 64'd0;
	mem_4[473] = 64'd0;
	mem_4[474] = 64'd0;
	mem_4[475] = 64'd0;
	mem_4[476] = 64'd0;
	mem_4[477] = 64'd0;
	mem_4[478] = 64'd0;
	mem_4[479] = 64'd0;
	mem_4[480] = 64'd0;
	mem_4[481] = 64'd0;
	mem_4[482] = 64'd0;
	mem_4[483] = 64'd0;
	mem_4[484] = 64'd0;
	mem_4[485] = 64'd0;
	mem_4[486] = 64'd0;
	mem_4[487] = 64'd0;
	mem_4[488] = 64'd0;
	mem_4[489] = 64'd0;
	mem_4[490] = 64'd0;
	mem_4[491] = 64'd0;
	mem_4[492] = 64'd0;
	mem_4[493] = 64'd0;
	mem_4[494] = 64'd0;
	mem_4[495] = 64'd0;
	mem_4[496] = 64'd0;
	mem_4[497] = 64'd0;
	mem_4[498] = 64'd0;
	mem_4[499] = 64'd0;
	mem_4[500] = 64'd0;
	mem_4[501] = 64'd0;
	mem_4[502] = 64'd0;
	mem_4[503] = 64'd0;
	mem_4[504] = 64'd0;
	mem_4[505] = 64'd0;
	mem_4[506] = 64'd0;
	mem_4[507] = 64'd0;
	mem_4[508] = 64'd0;
	mem_4[509] = 64'd0;
	mem_4[510] = 64'd0;
	mem_4[511] = 64'd0;
	mem_4[512] = 64'd0;
	mem_4[513] = 64'd0;
	mem_4[514] = 64'd0;
	mem_4[515] = 64'd0;
	mem_4[516] = 64'd0;
	mem_4[517] = 64'd0;
	mem_4[518] = 64'd0;
	mem_4[519] = 64'd0;
	mem_4[520] = 64'd0;
	mem_4[521] = 64'd0;
	mem_4[522] = 64'd0;
	mem_4[523] = 64'd0;
	mem_4[524] = 64'd0;
	mem_4[525] = 64'd0;
	mem_4[526] = 64'd0;
	mem_4[527] = 64'd0;
	mem_4[528] = 64'd0;
	mem_4[529] = 64'd0;
	mem_4[530] = 64'd0;
	mem_4[531] = 64'd0;
	mem_4[532] = 64'd0;
	mem_4[533] = 64'd0;
	mem_4[534] = 64'd0;
	mem_4[535] = 64'd0;
	mem_4[536] = 64'd0;
	mem_4[537] = 64'd0;
	mem_4[538] = 64'd0;
	mem_4[539] = 64'd0;
	mem_4[540] = 64'd0;
	mem_4[541] = 64'd0;
	mem_4[542] = 64'd0;
	mem_4[543] = 64'd0;
	mem_4[544] = 64'd0;
	mem_4[545] = 64'd0;
	mem_4[546] = 64'd0;
	mem_4[547] = 64'd0;
	mem_4[548] = 64'd0;
	mem_4[549] = 64'd0;
	mem_4[550] = 64'd0;
	mem_4[551] = 64'd0;
	mem_4[552] = 64'd0;
	mem_4[553] = 64'd0;
	mem_4[554] = 64'd0;
	mem_4[555] = 64'd0;
	mem_4[556] = 64'd0;
	mem_4[557] = 64'd0;
	mem_4[558] = 64'd0;
	mem_4[559] = 64'd0;
	mem_4[560] = 64'd0;
	mem_4[561] = 64'd0;
	mem_4[562] = 64'd0;
	mem_4[563] = 64'd0;
	mem_4[564] = 64'd0;
	mem_4[565] = 64'd0;
	mem_4[566] = 64'd0;
	mem_4[567] = 64'd0;
	mem_4[568] = 64'd0;
	mem_4[569] = 64'd0;
	mem_4[570] = 64'd0;
	mem_4[571] = 64'd0;
	mem_4[572] = 64'd0;
	mem_4[573] = 64'd0;
	mem_4[574] = 64'd0;
	mem_4[575] = 64'd0;
	mem_4[576] = 64'd0;
	mem_4[577] = 64'd0;
	mem_4[578] = 64'd0;
	mem_4[579] = 64'd0;
	mem_4[580] = 64'd0;
	mem_4[581] = 64'd0;
	mem_4[582] = 64'd0;
	mem_4[583] = 64'd0;
	mem_4[584] = 64'd0;
	mem_4[585] = 64'd0;
	mem_4[586] = 64'd0;
	mem_4[587] = 64'd0;
	mem_4[588] = 64'd0;
	mem_4[589] = 64'd0;
	mem_4[590] = 64'd0;
	mem_4[591] = 64'd0;
	mem_4[592] = 64'd0;
	mem_4[593] = 64'd0;
	mem_4[594] = 64'd0;
	mem_4[595] = 64'd0;
	mem_4[596] = 64'd0;
	mem_4[597] = 64'd0;
	mem_4[598] = 64'd0;
	mem_4[599] = 64'd0;
	mem_4[600] = 64'd0;
	mem_4[601] = 64'd0;
	mem_4[602] = 64'd0;
	mem_4[603] = 64'd0;
	mem_4[604] = 64'd0;
	mem_4[605] = 64'd0;
	mem_4[606] = 64'd0;
	mem_4[607] = 64'd0;
	mem_4[608] = 64'd0;
	mem_4[609] = 64'd0;
	mem_4[610] = 64'd0;
	mem_4[611] = 64'd0;
	mem_4[612] = 64'd0;
	mem_4[613] = 64'd0;
	mem_4[614] = 64'd0;
	mem_4[615] = 64'd0;
	mem_4[616] = 64'd0;
	mem_4[617] = 64'd0;
	mem_4[618] = 64'd0;
	mem_4[619] = 64'd0;
	mem_4[620] = 64'd0;
	mem_4[621] = 64'd0;
	mem_4[622] = 64'd0;
	mem_4[623] = 64'd0;
	mem_4[624] = 64'd0;
	mem_4[625] = 64'd0;
	mem_4[626] = 64'd0;
	mem_4[627] = 64'd0;
	mem_4[628] = 64'd0;
	mem_4[629] = 64'd0;
	mem_4[630] = 64'd0;
	mem_4[631] = 64'd0;
	mem_4[632] = 64'd0;
	mem_4[633] = 64'd0;
	mem_4[634] = 64'd0;
	mem_4[635] = 64'd0;
	mem_4[636] = 64'd0;
	mem_4[637] = 64'd0;
	mem_4[638] = 64'd0;
	mem_4[639] = 64'd0;
	mem_4[640] = 64'd0;
	mem_4[641] = 64'd0;
	mem_4[642] = 64'd0;
	mem_4[643] = 64'd0;
	mem_4[644] = 64'd0;
	mem_4[645] = 64'd0;
	mem_4[646] = 64'd0;
	mem_4[647] = 64'd0;
	mem_4[648] = 64'd0;
	mem_4[649] = 64'd0;
	mem_4[650] = 64'd0;
	mem_4[651] = 64'd0;
	mem_4[652] = 64'd0;
	mem_4[653] = 64'd0;
	mem_4[654] = 64'd0;
	mem_4[655] = 64'd0;
	mem_4[656] = 64'd0;
	mem_4[657] = 64'd0;
	mem_4[658] = 64'd0;
	mem_4[659] = 64'd0;
	mem_4[660] = 64'd0;
	mem_4[661] = 64'd0;
	mem_4[662] = 64'd0;
	mem_4[663] = 64'd0;
	mem_4[664] = 64'd0;
	mem_4[665] = 64'd0;
	mem_4[666] = 64'd0;
	mem_4[667] = 64'd0;
	mem_4[668] = 64'd0;
	mem_4[669] = 64'd0;
	mem_4[670] = 64'd0;
	mem_4[671] = 64'd0;
	mem_4[672] = 64'd0;
	mem_4[673] = 64'd0;
	mem_4[674] = 64'd0;
	mem_4[675] = 64'd0;
	mem_4[676] = 64'd0;
	mem_4[677] = 64'd0;
	mem_4[678] = 64'd0;
	mem_4[679] = 64'd0;
	mem_4[680] = 64'd0;
	mem_4[681] = 64'd0;
	mem_4[682] = 64'd0;
	mem_4[683] = 64'd0;
	mem_4[684] = 64'd0;
	mem_4[685] = 64'd0;
	mem_4[686] = 64'd0;
	mem_4[687] = 64'd0;
	mem_4[688] = 64'd0;
	mem_4[689] = 64'd0;
	mem_4[690] = 64'd0;
	mem_4[691] = 64'd0;
	mem_4[692] = 64'd0;
	mem_4[693] = 64'd0;
	mem_4[694] = 64'd0;
	mem_4[695] = 64'd0;
	mem_4[696] = 64'd0;
	mem_4[697] = 64'd0;
	mem_4[698] = 64'd0;
	mem_4[699] = 64'd0;
	mem_4[700] = 64'd0;
	mem_4[701] = 64'd0;
	mem_4[702] = 64'd0;
	mem_4[703] = 64'd0;
	mem_4[704] = 64'd0;
	mem_4[705] = 64'd0;
	mem_4[706] = 64'd0;
	mem_4[707] = 64'd0;
	mem_4[708] = 64'd0;
	mem_4[709] = 64'd0;
	mem_4[710] = 64'd0;
	mem_4[711] = 64'd0;
	mem_4[712] = 64'd0;
	mem_4[713] = 64'd0;
	mem_4[714] = 64'd0;
	mem_4[715] = 64'd0;
	mem_4[716] = 64'd0;
	mem_4[717] = 64'd0;
	mem_4[718] = 64'd0;
	mem_4[719] = 64'd0;
	mem_4[720] = 64'd0;
	mem_4[721] = 64'd0;
	mem_4[722] = 64'd0;
	mem_4[723] = 64'd0;
	mem_4[724] = 64'd0;
	mem_4[725] = 64'd0;
	mem_4[726] = 64'd0;
	mem_4[727] = 64'd0;
	mem_4[728] = 64'd0;
	mem_4[729] = 64'd0;
	mem_4[730] = 64'd0;
	mem_4[731] = 64'd0;
	mem_4[732] = 64'd0;
	mem_4[733] = 64'd0;
	mem_4[734] = 64'd0;
	mem_4[735] = 64'd0;
	mem_4[736] = 64'd0;
	mem_4[737] = 64'd0;
	mem_4[738] = 64'd0;
	mem_4[739] = 64'd0;
	mem_4[740] = 64'd0;
	mem_4[741] = 64'd0;
	mem_4[742] = 64'd0;
	mem_4[743] = 64'd0;
	mem_4[744] = 64'd0;
	mem_4[745] = 64'd0;
	mem_4[746] = 64'd0;
	mem_4[747] = 64'd0;
	mem_4[748] = 64'd0;
	mem_4[749] = 64'd0;
	mem_4[750] = 64'd0;
	mem_4[751] = 64'd0;
	mem_4[752] = 64'd0;
	mem_4[753] = 64'd0;
	mem_4[754] = 64'd0;
	mem_4[755] = 64'd0;
	mem_4[756] = 64'd0;
	mem_4[757] = 64'd0;
	mem_4[758] = 64'd0;
	mem_4[759] = 64'd0;
	mem_4[760] = 64'd0;
	mem_4[761] = 64'd0;
	mem_4[762] = 64'd0;
	mem_4[763] = 64'd0;
	mem_4[764] = 64'd0;
	mem_4[765] = 64'd0;
	mem_4[766] = 64'd0;
	mem_4[767] = 64'd0;
	mem_4[768] = 64'd0;
	mem_4[769] = 64'd0;
	mem_4[770] = 64'd0;
	mem_4[771] = 64'd0;
	mem_4[772] = 64'd0;
	mem_4[773] = 64'd0;
	mem_4[774] = 64'd0;
	mem_4[775] = 64'd0;
	mem_4[776] = 64'd0;
	mem_4[777] = 64'd0;
	mem_4[778] = 64'd0;
	mem_4[779] = 64'd0;
	mem_4[780] = 64'd0;
	mem_4[781] = 64'd0;
	mem_4[782] = 64'd0;
	mem_4[783] = 64'd0;
	mem_4[784] = 64'd0;
	mem_4[785] = 64'd0;
	mem_4[786] = 64'd0;
	mem_4[787] = 64'd0;
	mem_4[788] = 64'd0;
	mem_4[789] = 64'd0;
	mem_4[790] = 64'd0;
	mem_4[791] = 64'd0;
	mem_4[792] = 64'd0;
	mem_4[793] = 64'd0;
	mem_4[794] = 64'd0;
	mem_4[795] = 64'd0;
	mem_4[796] = 64'd0;
	mem_4[797] = 64'd0;
	mem_4[798] = 64'd0;
	mem_4[799] = 64'd0;
	mem_4[800] = 64'd0;
	mem_4[801] = 64'd0;
	mem_4[802] = 64'd0;
	mem_4[803] = 64'd0;
	mem_4[804] = 64'd0;
	mem_4[805] = 64'd0;
	mem_4[806] = 64'd0;
	mem_4[807] = 64'd0;
	mem_4[808] = 64'd0;
	mem_4[809] = 64'd0;
	mem_4[810] = 64'd0;
	mem_4[811] = 64'd0;
	mem_4[812] = 64'd0;
	mem_4[813] = 64'd0;
	mem_4[814] = 64'd0;
	mem_4[815] = 64'd0;
	mem_4[816] = 64'd0;
	mem_4[817] = 64'd0;
	mem_4[818] = 64'd0;
	mem_4[819] = 64'd0;
	mem_4[820] = 64'd0;
	mem_4[821] = 64'd0;
	mem_4[822] = 64'd0;
	mem_4[823] = 64'd0;
	mem_4[824] = 64'd0;
	mem_4[825] = 64'd0;
	mem_4[826] = 64'd0;
	mem_4[827] = 64'd0;
	mem_4[828] = 64'd0;
	mem_4[829] = 64'd0;
	mem_4[830] = 64'd0;
	mem_4[831] = 64'd0;
	mem_4[832] = 64'd0;
	mem_4[833] = 64'd0;
	mem_4[834] = 64'd0;
	mem_4[835] = 64'd0;
	mem_4[836] = 64'd0;
	mem_4[837] = 64'd0;
	mem_4[838] = 64'd0;
	mem_4[839] = 64'd0;
	mem_4[840] = 64'd0;
	mem_4[841] = 64'd0;
	mem_4[842] = 64'd0;
	mem_4[843] = 64'd0;
	mem_4[844] = 64'd0;
	mem_4[845] = 64'd0;
	mem_4[846] = 64'd0;
	mem_4[847] = 64'd0;
	mem_4[848] = 64'd0;
	mem_4[849] = 64'd0;
	mem_4[850] = 64'd0;
	mem_4[851] = 64'd0;
	mem_4[852] = 64'd0;
	mem_4[853] = 64'd0;
	mem_4[854] = 64'd0;
	mem_4[855] = 64'd0;
	mem_4[856] = 64'd0;
	mem_4[857] = 64'd0;
	mem_4[858] = 64'd0;
	mem_4[859] = 64'd0;
	mem_4[860] = 64'd0;
	mem_4[861] = 64'd0;
	mem_4[862] = 64'd0;
	mem_4[863] = 64'd0;
	mem_4[864] = 64'd0;
	mem_4[865] = 64'd0;
	mem_4[866] = 64'd0;
	mem_4[867] = 64'd0;
	mem_4[868] = 64'd0;
	mem_4[869] = 64'd0;
	mem_4[870] = 64'd0;
	mem_4[871] = 64'd0;
	mem_4[872] = 64'd0;
	mem_4[873] = 64'd0;
	mem_4[874] = 64'd0;
	mem_4[875] = 64'd0;
	mem_4[876] = 64'd0;
	mem_4[877] = 64'd0;
	mem_4[878] = 64'd0;
	mem_4[879] = 64'd0;
	mem_4[880] = 64'd0;
	mem_4[881] = 64'd0;
	mem_4[882] = 64'd0;
	mem_4[883] = 64'd0;
	mem_4[884] = 64'd0;
	mem_4[885] = 64'd0;
	mem_4[886] = 64'd0;
	mem_4[887] = 64'd0;
	mem_4[888] = 64'd0;
	mem_4[889] = 64'd0;
	mem_4[890] = 64'd0;
	mem_4[891] = 64'd0;
	mem_4[892] = 64'd0;
	mem_4[893] = 64'd0;
	mem_4[894] = 64'd0;
	mem_4[895] = 64'd0;
	mem_4[896] = 64'd0;
	mem_4[897] = 64'd0;
	mem_4[898] = 64'd0;
	mem_4[899] = 64'd0;
	mem_4[900] = 64'd0;
	mem_4[901] = 64'd0;
	mem_4[902] = 64'd0;
	mem_4[903] = 64'd0;
	mem_4[904] = 64'd0;
	mem_4[905] = 64'd0;
	mem_4[906] = 64'd0;
	mem_4[907] = 64'd0;
	mem_4[908] = 64'd0;
	mem_4[909] = 64'd0;
	mem_4[910] = 64'd0;
	mem_4[911] = 64'd0;
	mem_4[912] = 64'd0;
	mem_4[913] = 64'd0;
	mem_4[914] = 64'd0;
	mem_4[915] = 64'd0;
	mem_4[916] = 64'd0;
	mem_4[917] = 64'd0;
	mem_4[918] = 64'd0;
	mem_4[919] = 64'd0;
	mem_4[920] = 64'd0;
	mem_4[921] = 64'd0;
	mem_4[922] = 64'd0;
	mem_4[923] = 64'd0;
	mem_4[924] = 64'd0;
	mem_4[925] = 64'd0;
	mem_4[926] = 64'd0;
	mem_4[927] = 64'd0;
	mem_4[928] = 64'd0;
	mem_4[929] = 64'd0;
	mem_4[930] = 64'd0;
	mem_4[931] = 64'd0;
	mem_4[932] = 64'd0;
	mem_4[933] = 64'd0;
	mem_4[934] = 64'd0;
	mem_4[935] = 64'd0;
	mem_4[936] = 64'd0;
	mem_4[937] = 64'd0;
	mem_4[938] = 64'd0;
	mem_4[939] = 64'd0;
	mem_4[940] = 64'd0;
	mem_4[941] = 64'd0;
	mem_4[942] = 64'd0;
	mem_4[943] = 64'd0;
	mem_4[944] = 64'd0;
	mem_4[945] = 64'd0;
	mem_4[946] = 64'd0;
	mem_4[947] = 64'd0;
	mem_4[948] = 64'd0;
	mem_4[949] = 64'd0;
	mem_4[950] = 64'd0;
	mem_4[951] = 64'd0;
	mem_4[952] = 64'd0;
	mem_4[953] = 64'd0;
	mem_4[954] = 64'd0;
	mem_4[955] = 64'd0;
	mem_4[956] = 64'd0;
	mem_4[957] = 64'd0;
	mem_4[958] = 64'd0;
	mem_4[959] = 64'd0;
	mem_4[960] = 64'd0;
	mem_4[961] = 64'd0;
	mem_4[962] = 64'd0;
	mem_4[963] = 64'd0;
	mem_4[964] = 64'd0;
	mem_4[965] = 64'd0;
	mem_4[966] = 64'd0;
	mem_4[967] = 64'd0;
	mem_4[968] = 64'd0;
	mem_4[969] = 64'd0;
	mem_4[970] = 64'd0;
	mem_4[971] = 64'd0;
	mem_4[972] = 64'd0;
	mem_4[973] = 64'd0;
	mem_4[974] = 64'd0;
	mem_4[975] = 64'd0;
	mem_4[976] = 64'd0;
	mem_4[977] = 64'd0;
	mem_4[978] = 64'd0;
	mem_4[979] = 64'd0;
	mem_4[980] = 64'd0;
	mem_4[981] = 64'd0;
	mem_4[982] = 64'd0;
	mem_4[983] = 64'd0;
	mem_4[984] = 64'd0;
	mem_4[985] = 64'd0;
	mem_4[986] = 64'd0;
	mem_4[987] = 64'd0;
	mem_4[988] = 64'd0;
	mem_4[989] = 64'd0;
	mem_4[990] = 64'd0;
	mem_4[991] = 64'd0;
	mem_4[992] = 64'd0;
	mem_4[993] = 64'd0;
	mem_4[994] = 64'd0;
	mem_4[995] = 64'd0;
	mem_4[996] = 64'd0;
	mem_4[997] = 64'd0;
	mem_4[998] = 64'd0;
	mem_4[999] = 64'd0;
	mem_4[1000] = 64'd0;
	mem_4[1001] = 64'd0;
	mem_4[1002] = 64'd0;
	mem_4[1003] = 64'd0;
	mem_4[1004] = 64'd0;
	mem_4[1005] = 64'd0;
	mem_4[1006] = 64'd0;
	mem_4[1007] = 64'd0;
	mem_4[1008] = 64'd0;
	mem_4[1009] = 64'd0;
	mem_4[1010] = 64'd0;
	mem_4[1011] = 64'd0;
	mem_4[1012] = 64'd0;
	mem_4[1013] = 64'd0;
	mem_4[1014] = 64'd0;
	mem_4[1015] = 64'd0;
	mem_4[1016] = 64'd0;
	mem_4[1017] = 64'd0;
	mem_4[1018] = 64'd0;
	mem_4[1019] = 64'd0;
	mem_4[1020] = 64'd0;
	mem_4[1021] = 64'd0;
	mem_4[1022] = 64'd0;
	mem_4[1023] = 64'd0;
	mem_5[0] = 64'd0;
	mem_5[1] = 64'd0;
	mem_5[2] = 64'd0;
	mem_5[3] = 64'd0;
	mem_5[4] = 64'd0;
	mem_5[5] = 64'd0;
	mem_5[6] = 64'd0;
	mem_5[7] = 64'd0;
	mem_5[8] = 64'd0;
	mem_5[9] = 64'd0;
	mem_5[10] = 64'd0;
	mem_5[11] = 64'd0;
	mem_5[12] = 64'd0;
	mem_5[13] = 64'd0;
	mem_5[14] = 64'd0;
	mem_5[15] = 64'd0;
	mem_5[16] = 64'd0;
	mem_5[17] = 64'd0;
	mem_5[18] = 64'd0;
	mem_5[19] = 64'd0;
	mem_5[20] = 64'd0;
	mem_5[21] = 64'd0;
	mem_5[22] = 64'd0;
	mem_5[23] = 64'd0;
	mem_5[24] = 64'd0;
	mem_5[25] = 64'd0;
	mem_5[26] = 64'd0;
	mem_5[27] = 64'd0;
	mem_5[28] = 64'd0;
	mem_5[29] = 64'd0;
	mem_5[30] = 64'd0;
	mem_5[31] = 64'd0;
	mem_5[32] = 64'd0;
	mem_5[33] = 64'd0;
	mem_5[34] = 64'd0;
	mem_5[35] = 64'd0;
	mem_5[36] = 64'd0;
	mem_5[37] = 64'd0;
	mem_5[38] = 64'd0;
	mem_5[39] = 64'd0;
	mem_5[40] = 64'd0;
	mem_5[41] = 64'd0;
	mem_5[42] = 64'd0;
	mem_5[43] = 64'd0;
	mem_5[44] = 64'd0;
	mem_5[45] = 64'd0;
	mem_5[46] = 64'd0;
	mem_5[47] = 64'd0;
	mem_5[48] = 64'd0;
	mem_5[49] = 64'd0;
	mem_5[50] = 64'd0;
	mem_5[51] = 64'd0;
	mem_5[52] = 64'd0;
	mem_5[53] = 64'd0;
	mem_5[54] = 64'd0;
	mem_5[55] = 64'd0;
	mem_5[56] = 64'd0;
	mem_5[57] = 64'd0;
	mem_5[58] = 64'd0;
	mem_5[59] = 64'd0;
	mem_5[60] = 64'd0;
	mem_5[61] = 64'd0;
	mem_5[62] = 64'd0;
	mem_5[63] = 64'd0;
	mem_5[64] = 64'd0;
	mem_5[65] = 64'd0;
	mem_5[66] = 64'd0;
	mem_5[67] = 64'd0;
	mem_5[68] = 64'd0;
	mem_5[69] = 64'd0;
	mem_5[70] = 64'd0;
	mem_5[71] = 64'd0;
	mem_5[72] = 64'd0;
	mem_5[73] = 64'd0;
	mem_5[74] = 64'd0;
	mem_5[75] = 64'd0;
	mem_5[76] = 64'd0;
	mem_5[77] = 64'd0;
	mem_5[78] = 64'd0;
	mem_5[79] = 64'd0;
	mem_5[80] = 64'd0;
	mem_5[81] = 64'd0;
	mem_5[82] = 64'd0;
	mem_5[83] = 64'd0;
	mem_5[84] = 64'd0;
	mem_5[85] = 64'd0;
	mem_5[86] = 64'd0;
	mem_5[87] = 64'd0;
	mem_5[88] = 64'd0;
	mem_5[89] = 64'd0;
	mem_5[90] = 64'd0;
	mem_5[91] = 64'd0;
	mem_5[92] = 64'd0;
	mem_5[93] = 64'd0;
	mem_5[94] = 64'd0;
	mem_5[95] = 64'd0;
	mem_5[96] = 64'd0;
	mem_5[97] = 64'd0;
	mem_5[98] = 64'd0;
	mem_5[99] = 64'd0;
	mem_5[100] = 64'd0;
	mem_5[101] = 64'd0;
	mem_5[102] = 64'd0;
	mem_5[103] = 64'd0;
	mem_5[104] = 64'd0;
	mem_5[105] = 64'd0;
	mem_5[106] = 64'd0;
	mem_5[107] = 64'd0;
	mem_5[108] = 64'd0;
	mem_5[109] = 64'd0;
	mem_5[110] = 64'd0;
	mem_5[111] = 64'd0;
	mem_5[112] = 64'd0;
	mem_5[113] = 64'd0;
	mem_5[114] = 64'd0;
	mem_5[115] = 64'd0;
	mem_5[116] = 64'd0;
	mem_5[117] = 64'd0;
	mem_5[118] = 64'd0;
	mem_5[119] = 64'd0;
	mem_5[120] = 64'd0;
	mem_5[121] = 64'd0;
	mem_5[122] = 64'd0;
	mem_5[123] = 64'd0;
	mem_5[124] = 64'd0;
	mem_5[125] = 64'd0;
	mem_5[126] = 64'd0;
	mem_5[127] = 64'd0;
	mem_5[128] = 64'd0;
	mem_5[129] = 64'd0;
	mem_5[130] = 64'd0;
	mem_5[131] = 64'd0;
	mem_5[132] = 64'd0;
	mem_5[133] = 64'd0;
	mem_5[134] = 64'd0;
	mem_5[135] = 64'd0;
	mem_5[136] = 64'd0;
	mem_5[137] = 64'd0;
	mem_5[138] = 64'd0;
	mem_5[139] = 64'd0;
	mem_5[140] = 64'd0;
	mem_5[141] = 64'd0;
	mem_5[142] = 64'd0;
	mem_5[143] = 64'd0;
	mem_5[144] = 64'd0;
	mem_5[145] = 64'd0;
	mem_5[146] = 64'd0;
	mem_5[147] = 64'd0;
	mem_5[148] = 64'd0;
	mem_5[149] = 64'd0;
	mem_5[150] = 64'd0;
	mem_5[151] = 64'd0;
	mem_5[152] = 64'd0;
	mem_5[153] = 64'd0;
	mem_5[154] = 64'd0;
	mem_5[155] = 64'd0;
	mem_5[156] = 64'd0;
	mem_5[157] = 64'd0;
	mem_5[158] = 64'd0;
	mem_5[159] = 64'd0;
	mem_5[160] = 64'd0;
	mem_5[161] = 64'd0;
	mem_5[162] = 64'd0;
	mem_5[163] = 64'd0;
	mem_5[164] = 64'd0;
	mem_5[165] = 64'd0;
	mem_5[166] = 64'd0;
	mem_5[167] = 64'd0;
	mem_5[168] = 64'd0;
	mem_5[169] = 64'd0;
	mem_5[170] = 64'd0;
	mem_5[171] = 64'd0;
	mem_5[172] = 64'd0;
	mem_5[173] = 64'd0;
	mem_5[174] = 64'd0;
	mem_5[175] = 64'd0;
	mem_5[176] = 64'd0;
	mem_5[177] = 64'd0;
	mem_5[178] = 64'd0;
	mem_5[179] = 64'd0;
	mem_5[180] = 64'd0;
	mem_5[181] = 64'd0;
	mem_5[182] = 64'd0;
	mem_5[183] = 64'd0;
	mem_5[184] = 64'd0;
	mem_5[185] = 64'd0;
	mem_5[186] = 64'd0;
	mem_5[187] = 64'd0;
	mem_5[188] = 64'd0;
	mem_5[189] = 64'd0;
	mem_5[190] = 64'd0;
	mem_5[191] = 64'd0;
	mem_5[192] = 64'd0;
	mem_5[193] = 64'd0;
	mem_5[194] = 64'd0;
	mem_5[195] = 64'd0;
	mem_5[196] = 64'd0;
	mem_5[197] = 64'd0;
	mem_5[198] = 64'd0;
	mem_5[199] = 64'd0;
	mem_5[200] = 64'd0;
	mem_5[201] = 64'd0;
	mem_5[202] = 64'd0;
	mem_5[203] = 64'd0;
	mem_5[204] = 64'd0;
	mem_5[205] = 64'd0;
	mem_5[206] = 64'd0;
	mem_5[207] = 64'd0;
	mem_5[208] = 64'd0;
	mem_5[209] = 64'd0;
	mem_5[210] = 64'd0;
	mem_5[211] = 64'd0;
	mem_5[212] = 64'd0;
	mem_5[213] = 64'd0;
	mem_5[214] = 64'd0;
	mem_5[215] = 64'd0;
	mem_5[216] = 64'd0;
	mem_5[217] = 64'd0;
	mem_5[218] = 64'd0;
	mem_5[219] = 64'd0;
	mem_5[220] = 64'd0;
	mem_5[221] = 64'd0;
	mem_5[222] = 64'd0;
	mem_5[223] = 64'd0;
	mem_5[224] = 64'd0;
	mem_5[225] = 64'd0;
	mem_5[226] = 64'd0;
	mem_5[227] = 64'd0;
	mem_5[228] = 64'd0;
	mem_5[229] = 64'd0;
	mem_5[230] = 64'd0;
	mem_5[231] = 64'd0;
	mem_5[232] = 64'd0;
	mem_5[233] = 64'd0;
	mem_5[234] = 64'd0;
	mem_5[235] = 64'd0;
	mem_5[236] = 64'd0;
	mem_5[237] = 64'd0;
	mem_5[238] = 64'd0;
	mem_5[239] = 64'd0;
	mem_5[240] = 64'd0;
	mem_5[241] = 64'd0;
	mem_5[242] = 64'd0;
	mem_5[243] = 64'd0;
	mem_5[244] = 64'd0;
	mem_5[245] = 64'd0;
	mem_5[246] = 64'd0;
	mem_5[247] = 64'd0;
	mem_5[248] = 64'd0;
	mem_5[249] = 64'd0;
	mem_5[250] = 64'd0;
	mem_5[251] = 64'd0;
	mem_5[252] = 64'd0;
	mem_5[253] = 64'd0;
	mem_5[254] = 64'd0;
	mem_5[255] = 64'd0;
	mem_5[256] = 64'd0;
	mem_5[257] = 64'd0;
	mem_5[258] = 64'd0;
	mem_5[259] = 64'd0;
	mem_5[260] = 64'd0;
	mem_5[261] = 64'd0;
	mem_5[262] = 64'd0;
	mem_5[263] = 64'd0;
	mem_5[264] = 64'd0;
	mem_5[265] = 64'd0;
	mem_5[266] = 64'd0;
	mem_5[267] = 64'd0;
	mem_5[268] = 64'd0;
	mem_5[269] = 64'd0;
	mem_5[270] = 64'd0;
	mem_5[271] = 64'd0;
	mem_5[272] = 64'd0;
	mem_5[273] = 64'd0;
	mem_5[274] = 64'd0;
	mem_5[275] = 64'd0;
	mem_5[276] = 64'd0;
	mem_5[277] = 64'd0;
	mem_5[278] = 64'd0;
	mem_5[279] = 64'd0;
	mem_5[280] = 64'd0;
	mem_5[281] = 64'd0;
	mem_5[282] = 64'd0;
	mem_5[283] = 64'd0;
	mem_5[284] = 64'd0;
	mem_5[285] = 64'd0;
	mem_5[286] = 64'd0;
	mem_5[287] = 64'd0;
	mem_5[288] = 64'd0;
	mem_5[289] = 64'd0;
	mem_5[290] = 64'd0;
	mem_5[291] = 64'd0;
	mem_5[292] = 64'd0;
	mem_5[293] = 64'd0;
	mem_5[294] = 64'd0;
	mem_5[295] = 64'd0;
	mem_5[296] = 64'd0;
	mem_5[297] = 64'd0;
	mem_5[298] = 64'd0;
	mem_5[299] = 64'd0;
	mem_5[300] = 64'd0;
	mem_5[301] = 64'd0;
	mem_5[302] = 64'd0;
	mem_5[303] = 64'd0;
	mem_5[304] = 64'd0;
	mem_5[305] = 64'd0;
	mem_5[306] = 64'd0;
	mem_5[307] = 64'd0;
	mem_5[308] = 64'd0;
	mem_5[309] = 64'd0;
	mem_5[310] = 64'd0;
	mem_5[311] = 64'd0;
	mem_5[312] = 64'd0;
	mem_5[313] = 64'd0;
	mem_5[314] = 64'd0;
	mem_5[315] = 64'd0;
	mem_5[316] = 64'd0;
	mem_5[317] = 64'd0;
	mem_5[318] = 64'd0;
	mem_5[319] = 64'd0;
	mem_5[320] = 64'd0;
	mem_5[321] = 64'd0;
	mem_5[322] = 64'd0;
	mem_5[323] = 64'd0;
	mem_5[324] = 64'd0;
	mem_5[325] = 64'd0;
	mem_5[326] = 64'd0;
	mem_5[327] = 64'd0;
	mem_5[328] = 64'd0;
	mem_5[329] = 64'd0;
	mem_5[330] = 64'd0;
	mem_5[331] = 64'd0;
	mem_5[332] = 64'd0;
	mem_5[333] = 64'd0;
	mem_5[334] = 64'd0;
	mem_5[335] = 64'd0;
	mem_5[336] = 64'd0;
	mem_5[337] = 64'd0;
	mem_5[338] = 64'd0;
	mem_5[339] = 64'd0;
	mem_5[340] = 64'd0;
	mem_5[341] = 64'd0;
	mem_5[342] = 64'd0;
	mem_5[343] = 64'd0;
	mem_5[344] = 64'd0;
	mem_5[345] = 64'd0;
	mem_5[346] = 64'd0;
	mem_5[347] = 64'd0;
	mem_5[348] = 64'd0;
	mem_5[349] = 64'd0;
	mem_5[350] = 64'd0;
	mem_5[351] = 64'd0;
	mem_5[352] = 64'd0;
	mem_5[353] = 64'd0;
	mem_5[354] = 64'd0;
	mem_5[355] = 64'd0;
	mem_5[356] = 64'd0;
	mem_5[357] = 64'd0;
	mem_5[358] = 64'd0;
	mem_5[359] = 64'd0;
	mem_5[360] = 64'd0;
	mem_5[361] = 64'd0;
	mem_5[362] = 64'd0;
	mem_5[363] = 64'd0;
	mem_5[364] = 64'd0;
	mem_5[365] = 64'd0;
	mem_5[366] = 64'd0;
	mem_5[367] = 64'd0;
	mem_5[368] = 64'd0;
	mem_5[369] = 64'd0;
	mem_5[370] = 64'd0;
	mem_5[371] = 64'd0;
	mem_5[372] = 64'd0;
	mem_5[373] = 64'd0;
	mem_5[374] = 64'd0;
	mem_5[375] = 64'd0;
	mem_5[376] = 64'd0;
	mem_5[377] = 64'd0;
	mem_5[378] = 64'd0;
	mem_5[379] = 64'd0;
	mem_5[380] = 64'd0;
	mem_5[381] = 64'd0;
	mem_5[382] = 64'd0;
	mem_5[383] = 64'd0;
	mem_5[384] = 64'd0;
	mem_5[385] = 64'd0;
	mem_5[386] = 64'd0;
	mem_5[387] = 64'd0;
	mem_5[388] = 64'd0;
	mem_5[389] = 64'd0;
	mem_5[390] = 64'd0;
	mem_5[391] = 64'd0;
	mem_5[392] = 64'd0;
	mem_5[393] = 64'd0;
	mem_5[394] = 64'd0;
	mem_5[395] = 64'd0;
	mem_5[396] = 64'd0;
	mem_5[397] = 64'd0;
	mem_5[398] = 64'd0;
	mem_5[399] = 64'd0;
	mem_5[400] = 64'd0;
	mem_5[401] = 64'd0;
	mem_5[402] = 64'd0;
	mem_5[403] = 64'd0;
	mem_5[404] = 64'd0;
	mem_5[405] = 64'd0;
	mem_5[406] = 64'd0;
	mem_5[407] = 64'd0;
	mem_5[408] = 64'd0;
	mem_5[409] = 64'd0;
	mem_5[410] = 64'd0;
	mem_5[411] = 64'd0;
	mem_5[412] = 64'd0;
	mem_5[413] = 64'd0;
	mem_5[414] = 64'd0;
	mem_5[415] = 64'd0;
	mem_5[416] = 64'd0;
	mem_5[417] = 64'd0;
	mem_5[418] = 64'd0;
	mem_5[419] = 64'd0;
	mem_5[420] = 64'd0;
	mem_5[421] = 64'd0;
	mem_5[422] = 64'd0;
	mem_5[423] = 64'd0;
	mem_5[424] = 64'd0;
	mem_5[425] = 64'd0;
	mem_5[426] = 64'd0;
	mem_5[427] = 64'd0;
	mem_5[428] = 64'd0;
	mem_5[429] = 64'd0;
	mem_5[430] = 64'd0;
	mem_5[431] = 64'd0;
	mem_5[432] = 64'd0;
	mem_5[433] = 64'd0;
	mem_5[434] = 64'd0;
	mem_5[435] = 64'd0;
	mem_5[436] = 64'd0;
	mem_5[437] = 64'd0;
	mem_5[438] = 64'd0;
	mem_5[439] = 64'd0;
	mem_5[440] = 64'd0;
	mem_5[441] = 64'd0;
	mem_5[442] = 64'd0;
	mem_5[443] = 64'd0;
	mem_5[444] = 64'd0;
	mem_5[445] = 64'd0;
	mem_5[446] = 64'd0;
	mem_5[447] = 64'd0;
	mem_5[448] = 64'd0;
	mem_5[449] = 64'd0;
	mem_5[450] = 64'd0;
	mem_5[451] = 64'd0;
	mem_5[452] = 64'd0;
	mem_5[453] = 64'd0;
	mem_5[454] = 64'd0;
	mem_5[455] = 64'd0;
	mem_5[456] = 64'd0;
	mem_5[457] = 64'd0;
	mem_5[458] = 64'd0;
	mem_5[459] = 64'd0;
	mem_5[460] = 64'd0;
	mem_5[461] = 64'd0;
	mem_5[462] = 64'd0;
	mem_5[463] = 64'd0;
	mem_5[464] = 64'd0;
	mem_5[465] = 64'd0;
	mem_5[466] = 64'd0;
	mem_5[467] = 64'd0;
	mem_5[468] = 64'd0;
	mem_5[469] = 64'd0;
	mem_5[470] = 64'd0;
	mem_5[471] = 64'd0;
	mem_5[472] = 64'd0;
	mem_5[473] = 64'd0;
	mem_5[474] = 64'd0;
	mem_5[475] = 64'd0;
	mem_5[476] = 64'd0;
	mem_5[477] = 64'd0;
	mem_5[478] = 64'd0;
	mem_5[479] = 64'd0;
	mem_5[480] = 64'd0;
	mem_5[481] = 64'd0;
	mem_5[482] = 64'd0;
	mem_5[483] = 64'd0;
	mem_5[484] = 64'd0;
	mem_5[485] = 64'd0;
	mem_5[486] = 64'd0;
	mem_5[487] = 64'd0;
	mem_5[488] = 64'd0;
	mem_5[489] = 64'd0;
	mem_5[490] = 64'd0;
	mem_5[491] = 64'd0;
	mem_5[492] = 64'd0;
	mem_5[493] = 64'd0;
	mem_5[494] = 64'd0;
	mem_5[495] = 64'd0;
	mem_5[496] = 64'd0;
	mem_5[497] = 64'd0;
	mem_5[498] = 64'd0;
	mem_5[499] = 64'd0;
	mem_5[500] = 64'd0;
	mem_5[501] = 64'd0;
	mem_5[502] = 64'd0;
	mem_5[503] = 64'd0;
	mem_5[504] = 64'd0;
	mem_5[505] = 64'd0;
	mem_5[506] = 64'd0;
	mem_5[507] = 64'd0;
	mem_5[508] = 64'd0;
	mem_5[509] = 64'd0;
	mem_5[510] = 64'd0;
	mem_5[511] = 64'd0;
	mem_5[512] = 64'd0;
	mem_5[513] = 64'd0;
	mem_5[514] = 64'd0;
	mem_5[515] = 64'd0;
	mem_5[516] = 64'd0;
	mem_5[517] = 64'd0;
	mem_5[518] = 64'd0;
	mem_5[519] = 64'd0;
	mem_5[520] = 64'd0;
	mem_5[521] = 64'd0;
	mem_5[522] = 64'd0;
	mem_5[523] = 64'd0;
	mem_5[524] = 64'd0;
	mem_5[525] = 64'd0;
	mem_5[526] = 64'd0;
	mem_5[527] = 64'd0;
	mem_5[528] = 64'd0;
	mem_5[529] = 64'd0;
	mem_5[530] = 64'd0;
	mem_5[531] = 64'd0;
	mem_5[532] = 64'd0;
	mem_5[533] = 64'd0;
	mem_5[534] = 64'd0;
	mem_5[535] = 64'd0;
	mem_5[536] = 64'd0;
	mem_5[537] = 64'd0;
	mem_5[538] = 64'd0;
	mem_5[539] = 64'd0;
	mem_5[540] = 64'd0;
	mem_5[541] = 64'd0;
	mem_5[542] = 64'd0;
	mem_5[543] = 64'd0;
	mem_5[544] = 64'd0;
	mem_5[545] = 64'd0;
	mem_5[546] = 64'd0;
	mem_5[547] = 64'd0;
	mem_5[548] = 64'd0;
	mem_5[549] = 64'd0;
	mem_5[550] = 64'd0;
	mem_5[551] = 64'd0;
	mem_5[552] = 64'd0;
	mem_5[553] = 64'd0;
	mem_5[554] = 64'd0;
	mem_5[555] = 64'd0;
	mem_5[556] = 64'd0;
	mem_5[557] = 64'd0;
	mem_5[558] = 64'd0;
	mem_5[559] = 64'd0;
	mem_5[560] = 64'd0;
	mem_5[561] = 64'd0;
	mem_5[562] = 64'd0;
	mem_5[563] = 64'd0;
	mem_5[564] = 64'd0;
	mem_5[565] = 64'd0;
	mem_5[566] = 64'd0;
	mem_5[567] = 64'd0;
	mem_5[568] = 64'd0;
	mem_5[569] = 64'd0;
	mem_5[570] = 64'd0;
	mem_5[571] = 64'd0;
	mem_5[572] = 64'd0;
	mem_5[573] = 64'd0;
	mem_5[574] = 64'd0;
	mem_5[575] = 64'd0;
	mem_5[576] = 64'd0;
	mem_5[577] = 64'd0;
	mem_5[578] = 64'd0;
	mem_5[579] = 64'd0;
	mem_5[580] = 64'd0;
	mem_5[581] = 64'd0;
	mem_5[582] = 64'd0;
	mem_5[583] = 64'd0;
	mem_5[584] = 64'd0;
	mem_5[585] = 64'd0;
	mem_5[586] = 64'd0;
	mem_5[587] = 64'd0;
	mem_5[588] = 64'd0;
	mem_5[589] = 64'd0;
	mem_5[590] = 64'd0;
	mem_5[591] = 64'd0;
	mem_5[592] = 64'd0;
	mem_5[593] = 64'd0;
	mem_5[594] = 64'd0;
	mem_5[595] = 64'd0;
	mem_5[596] = 64'd0;
	mem_5[597] = 64'd0;
	mem_5[598] = 64'd0;
	mem_5[599] = 64'd0;
	mem_5[600] = 64'd0;
	mem_5[601] = 64'd0;
	mem_5[602] = 64'd0;
	mem_5[603] = 64'd0;
	mem_5[604] = 64'd0;
	mem_5[605] = 64'd0;
	mem_5[606] = 64'd0;
	mem_5[607] = 64'd0;
	mem_5[608] = 64'd0;
	mem_5[609] = 64'd0;
	mem_5[610] = 64'd0;
	mem_5[611] = 64'd0;
	mem_5[612] = 64'd0;
	mem_5[613] = 64'd0;
	mem_5[614] = 64'd0;
	mem_5[615] = 64'd0;
	mem_5[616] = 64'd0;
	mem_5[617] = 64'd0;
	mem_5[618] = 64'd0;
	mem_5[619] = 64'd0;
	mem_5[620] = 64'd0;
	mem_5[621] = 64'd0;
	mem_5[622] = 64'd0;
	mem_5[623] = 64'd0;
	mem_5[624] = 64'd0;
	mem_5[625] = 64'd0;
	mem_5[626] = 64'd0;
	mem_5[627] = 64'd0;
	mem_5[628] = 64'd0;
	mem_5[629] = 64'd0;
	mem_5[630] = 64'd0;
	mem_5[631] = 64'd0;
	mem_5[632] = 64'd0;
	mem_5[633] = 64'd0;
	mem_5[634] = 64'd0;
	mem_5[635] = 64'd0;
	mem_5[636] = 64'd0;
	mem_5[637] = 64'd0;
	mem_5[638] = 64'd0;
	mem_5[639] = 64'd0;
	mem_5[640] = 64'd0;
	mem_5[641] = 64'd0;
	mem_5[642] = 64'd0;
	mem_5[643] = 64'd0;
	mem_5[644] = 64'd0;
	mem_5[645] = 64'd0;
	mem_5[646] = 64'd0;
	mem_5[647] = 64'd0;
	mem_5[648] = 64'd0;
	mem_5[649] = 64'd0;
	mem_5[650] = 64'd0;
	mem_5[651] = 64'd0;
	mem_5[652] = 64'd0;
	mem_5[653] = 64'd0;
	mem_5[654] = 64'd0;
	mem_5[655] = 64'd0;
	mem_5[656] = 64'd0;
	mem_5[657] = 64'd0;
	mem_5[658] = 64'd0;
	mem_5[659] = 64'd0;
	mem_5[660] = 64'd0;
	mem_5[661] = 64'd0;
	mem_5[662] = 64'd0;
	mem_5[663] = 64'd0;
	mem_5[664] = 64'd0;
	mem_5[665] = 64'd0;
	mem_5[666] = 64'd0;
	mem_5[667] = 64'd0;
	mem_5[668] = 64'd0;
	mem_5[669] = 64'd0;
	mem_5[670] = 64'd0;
	mem_5[671] = 64'd0;
	mem_5[672] = 64'd0;
	mem_5[673] = 64'd0;
	mem_5[674] = 64'd0;
	mem_5[675] = 64'd0;
	mem_5[676] = 64'd0;
	mem_5[677] = 64'd0;
	mem_5[678] = 64'd0;
	mem_5[679] = 64'd0;
	mem_5[680] = 64'd0;
	mem_5[681] = 64'd0;
	mem_5[682] = 64'd0;
	mem_5[683] = 64'd0;
	mem_5[684] = 64'd0;
	mem_5[685] = 64'd0;
	mem_5[686] = 64'd0;
	mem_5[687] = 64'd0;
	mem_5[688] = 64'd0;
	mem_5[689] = 64'd0;
	mem_5[690] = 64'd0;
	mem_5[691] = 64'd0;
	mem_5[692] = 64'd0;
	mem_5[693] = 64'd0;
	mem_5[694] = 64'd0;
	mem_5[695] = 64'd0;
	mem_5[696] = 64'd0;
	mem_5[697] = 64'd0;
	mem_5[698] = 64'd0;
	mem_5[699] = 64'd0;
	mem_5[700] = 64'd0;
	mem_5[701] = 64'd0;
	mem_5[702] = 64'd0;
	mem_5[703] = 64'd0;
	mem_5[704] = 64'd0;
	mem_5[705] = 64'd0;
	mem_5[706] = 64'd0;
	mem_5[707] = 64'd0;
	mem_5[708] = 64'd0;
	mem_5[709] = 64'd0;
	mem_5[710] = 64'd0;
	mem_5[711] = 64'd0;
	mem_5[712] = 64'd0;
	mem_5[713] = 64'd0;
	mem_5[714] = 64'd0;
	mem_5[715] = 64'd0;
	mem_5[716] = 64'd0;
	mem_5[717] = 64'd0;
	mem_5[718] = 64'd0;
	mem_5[719] = 64'd0;
	mem_5[720] = 64'd0;
	mem_5[721] = 64'd0;
	mem_5[722] = 64'd0;
	mem_5[723] = 64'd0;
	mem_5[724] = 64'd0;
	mem_5[725] = 64'd0;
	mem_5[726] = 64'd0;
	mem_5[727] = 64'd0;
	mem_5[728] = 64'd0;
	mem_5[729] = 64'd0;
	mem_5[730] = 64'd0;
	mem_5[731] = 64'd0;
	mem_5[732] = 64'd0;
	mem_5[733] = 64'd0;
	mem_5[734] = 64'd0;
	mem_5[735] = 64'd0;
	mem_5[736] = 64'd0;
	mem_5[737] = 64'd0;
	mem_5[738] = 64'd0;
	mem_5[739] = 64'd0;
	mem_5[740] = 64'd0;
	mem_5[741] = 64'd0;
	mem_5[742] = 64'd0;
	mem_5[743] = 64'd0;
	mem_5[744] = 64'd0;
	mem_5[745] = 64'd0;
	mem_5[746] = 64'd0;
	mem_5[747] = 64'd0;
	mem_5[748] = 64'd0;
	mem_5[749] = 64'd0;
	mem_5[750] = 64'd0;
	mem_5[751] = 64'd0;
	mem_5[752] = 64'd0;
	mem_5[753] = 64'd0;
	mem_5[754] = 64'd0;
	mem_5[755] = 64'd0;
	mem_5[756] = 64'd0;
	mem_5[757] = 64'd0;
	mem_5[758] = 64'd0;
	mem_5[759] = 64'd0;
	mem_5[760] = 64'd0;
	mem_5[761] = 64'd0;
	mem_5[762] = 64'd0;
	mem_5[763] = 64'd0;
	mem_5[764] = 64'd0;
	mem_5[765] = 64'd0;
	mem_5[766] = 64'd0;
	mem_5[767] = 64'd0;
	mem_5[768] = 64'd0;
	mem_5[769] = 64'd0;
	mem_5[770] = 64'd0;
	mem_5[771] = 64'd0;
	mem_5[772] = 64'd0;
	mem_5[773] = 64'd0;
	mem_5[774] = 64'd0;
	mem_5[775] = 64'd0;
	mem_5[776] = 64'd0;
	mem_5[777] = 64'd0;
	mem_5[778] = 64'd0;
	mem_5[779] = 64'd0;
	mem_5[780] = 64'd0;
	mem_5[781] = 64'd0;
	mem_5[782] = 64'd0;
	mem_5[783] = 64'd0;
	mem_5[784] = 64'd0;
	mem_5[785] = 64'd0;
	mem_5[786] = 64'd0;
	mem_5[787] = 64'd0;
	mem_5[788] = 64'd0;
	mem_5[789] = 64'd0;
	mem_5[790] = 64'd0;
	mem_5[791] = 64'd0;
	mem_5[792] = 64'd0;
	mem_5[793] = 64'd0;
	mem_5[794] = 64'd0;
	mem_5[795] = 64'd0;
	mem_5[796] = 64'd0;
	mem_5[797] = 64'd0;
	mem_5[798] = 64'd0;
	mem_5[799] = 64'd0;
	mem_5[800] = 64'd0;
	mem_5[801] = 64'd0;
	mem_5[802] = 64'd0;
	mem_5[803] = 64'd0;
	mem_5[804] = 64'd0;
	mem_5[805] = 64'd0;
	mem_5[806] = 64'd0;
	mem_5[807] = 64'd0;
	mem_5[808] = 64'd0;
	mem_5[809] = 64'd0;
	mem_5[810] = 64'd0;
	mem_5[811] = 64'd0;
	mem_5[812] = 64'd0;
	mem_5[813] = 64'd0;
	mem_5[814] = 64'd0;
	mem_5[815] = 64'd0;
	mem_5[816] = 64'd0;
	mem_5[817] = 64'd0;
	mem_5[818] = 64'd0;
	mem_5[819] = 64'd0;
	mem_5[820] = 64'd0;
	mem_5[821] = 64'd0;
	mem_5[822] = 64'd0;
	mem_5[823] = 64'd0;
	mem_5[824] = 64'd0;
	mem_5[825] = 64'd0;
	mem_5[826] = 64'd0;
	mem_5[827] = 64'd0;
	mem_5[828] = 64'd0;
	mem_5[829] = 64'd0;
	mem_5[830] = 64'd0;
	mem_5[831] = 64'd0;
	mem_5[832] = 64'd0;
	mem_5[833] = 64'd0;
	mem_5[834] = 64'd0;
	mem_5[835] = 64'd0;
	mem_5[836] = 64'd0;
	mem_5[837] = 64'd0;
	mem_5[838] = 64'd0;
	mem_5[839] = 64'd0;
	mem_5[840] = 64'd0;
	mem_5[841] = 64'd0;
	mem_5[842] = 64'd0;
	mem_5[843] = 64'd0;
	mem_5[844] = 64'd0;
	mem_5[845] = 64'd0;
	mem_5[846] = 64'd0;
	mem_5[847] = 64'd0;
	mem_5[848] = 64'd0;
	mem_5[849] = 64'd0;
	mem_5[850] = 64'd0;
	mem_5[851] = 64'd0;
	mem_5[852] = 64'd0;
	mem_5[853] = 64'd0;
	mem_5[854] = 64'd0;
	mem_5[855] = 64'd0;
	mem_5[856] = 64'd0;
	mem_5[857] = 64'd0;
	mem_5[858] = 64'd0;
	mem_5[859] = 64'd0;
	mem_5[860] = 64'd0;
	mem_5[861] = 64'd0;
	mem_5[862] = 64'd0;
	mem_5[863] = 64'd0;
	mem_5[864] = 64'd0;
	mem_5[865] = 64'd0;
	mem_5[866] = 64'd0;
	mem_5[867] = 64'd0;
	mem_5[868] = 64'd0;
	mem_5[869] = 64'd0;
	mem_5[870] = 64'd0;
	mem_5[871] = 64'd0;
	mem_5[872] = 64'd0;
	mem_5[873] = 64'd0;
	mem_5[874] = 64'd0;
	mem_5[875] = 64'd0;
	mem_5[876] = 64'd0;
	mem_5[877] = 64'd0;
	mem_5[878] = 64'd0;
	mem_5[879] = 64'd0;
	mem_5[880] = 64'd0;
	mem_5[881] = 64'd0;
	mem_5[882] = 64'd0;
	mem_5[883] = 64'd0;
	mem_5[884] = 64'd0;
	mem_5[885] = 64'd0;
	mem_5[886] = 64'd0;
	mem_5[887] = 64'd0;
	mem_5[888] = 64'd0;
	mem_5[889] = 64'd0;
	mem_5[890] = 64'd0;
	mem_5[891] = 64'd0;
	mem_5[892] = 64'd0;
	mem_5[893] = 64'd0;
	mem_5[894] = 64'd0;
	mem_5[895] = 64'd0;
	mem_5[896] = 64'd0;
	mem_5[897] = 64'd0;
	mem_5[898] = 64'd0;
	mem_5[899] = 64'd0;
	mem_5[900] = 64'd0;
	mem_5[901] = 64'd0;
	mem_5[902] = 64'd0;
	mem_5[903] = 64'd0;
	mem_5[904] = 64'd0;
	mem_5[905] = 64'd0;
	mem_5[906] = 64'd0;
	mem_5[907] = 64'd0;
	mem_5[908] = 64'd0;
	mem_5[909] = 64'd0;
	mem_5[910] = 64'd0;
	mem_5[911] = 64'd0;
	mem_5[912] = 64'd0;
	mem_5[913] = 64'd0;
	mem_5[914] = 64'd0;
	mem_5[915] = 64'd0;
	mem_5[916] = 64'd0;
	mem_5[917] = 64'd0;
	mem_5[918] = 64'd0;
	mem_5[919] = 64'd0;
	mem_5[920] = 64'd0;
	mem_5[921] = 64'd0;
	mem_5[922] = 64'd0;
	mem_5[923] = 64'd0;
	mem_5[924] = 64'd0;
	mem_5[925] = 64'd0;
	mem_5[926] = 64'd0;
	mem_5[927] = 64'd0;
	mem_5[928] = 64'd0;
	mem_5[929] = 64'd0;
	mem_5[930] = 64'd0;
	mem_5[931] = 64'd0;
	mem_5[932] = 64'd0;
	mem_5[933] = 64'd0;
	mem_5[934] = 64'd0;
	mem_5[935] = 64'd0;
	mem_5[936] = 64'd0;
	mem_5[937] = 64'd0;
	mem_5[938] = 64'd0;
	mem_5[939] = 64'd0;
	mem_5[940] = 64'd0;
	mem_5[941] = 64'd0;
	mem_5[942] = 64'd0;
	mem_5[943] = 64'd0;
	mem_5[944] = 64'd0;
	mem_5[945] = 64'd0;
	mem_5[946] = 64'd0;
	mem_5[947] = 64'd0;
	mem_5[948] = 64'd0;
	mem_5[949] = 64'd0;
	mem_5[950] = 64'd0;
	mem_5[951] = 64'd0;
	mem_5[952] = 64'd0;
	mem_5[953] = 64'd0;
	mem_5[954] = 64'd0;
	mem_5[955] = 64'd0;
	mem_5[956] = 64'd0;
	mem_5[957] = 64'd0;
	mem_5[958] = 64'd0;
	mem_5[959] = 64'd0;
	mem_5[960] = 64'd0;
	mem_5[961] = 64'd0;
	mem_5[962] = 64'd0;
	mem_5[963] = 64'd0;
	mem_5[964] = 64'd0;
	mem_5[965] = 64'd0;
	mem_5[966] = 64'd0;
	mem_5[967] = 64'd0;
	mem_5[968] = 64'd0;
	mem_5[969] = 64'd0;
	mem_5[970] = 64'd0;
	mem_5[971] = 64'd0;
	mem_5[972] = 64'd0;
	mem_5[973] = 64'd0;
	mem_5[974] = 64'd0;
	mem_5[975] = 64'd0;
	mem_5[976] = 64'd0;
	mem_5[977] = 64'd0;
	mem_5[978] = 64'd0;
	mem_5[979] = 64'd0;
	mem_5[980] = 64'd0;
	mem_5[981] = 64'd0;
	mem_5[982] = 64'd0;
	mem_5[983] = 64'd0;
	mem_5[984] = 64'd0;
	mem_5[985] = 64'd0;
	mem_5[986] = 64'd0;
	mem_5[987] = 64'd0;
	mem_5[988] = 64'd0;
	mem_5[989] = 64'd0;
	mem_5[990] = 64'd0;
	mem_5[991] = 64'd0;
	mem_5[992] = 64'd0;
	mem_5[993] = 64'd0;
	mem_5[994] = 64'd0;
	mem_5[995] = 64'd0;
	mem_5[996] = 64'd0;
	mem_5[997] = 64'd0;
	mem_5[998] = 64'd0;
	mem_5[999] = 64'd0;
	mem_5[1000] = 64'd0;
	mem_5[1001] = 64'd0;
	mem_5[1002] = 64'd0;
	mem_5[1003] = 64'd0;
	mem_5[1004] = 64'd0;
	mem_5[1005] = 64'd0;
	mem_5[1006] = 64'd0;
	mem_5[1007] = 64'd0;
	mem_5[1008] = 64'd0;
	mem_5[1009] = 64'd0;
	mem_5[1010] = 64'd0;
	mem_5[1011] = 64'd0;
	mem_5[1012] = 64'd0;
	mem_5[1013] = 64'd0;
	mem_5[1014] = 64'd0;
	mem_5[1015] = 64'd0;
	mem_5[1016] = 64'd0;
	mem_5[1017] = 64'd0;
	mem_5[1018] = 64'd0;
	mem_5[1019] = 64'd0;
	mem_5[1020] = 64'd0;
	mem_5[1021] = 64'd0;
	mem_5[1022] = 64'd0;
	mem_5[1023] = 64'd0;
	mem_6[0] = 64'd0;
	mem_6[1] = 64'd0;
	mem_6[2] = 64'd0;
	mem_6[3] = 64'd0;
	mem_6[4] = 64'd0;
	mem_6[5] = 64'd0;
	mem_6[6] = 64'd0;
	mem_6[7] = 64'd0;
	mem_6[8] = 64'd0;
	mem_6[9] = 64'd0;
	mem_6[10] = 64'd0;
	mem_6[11] = 64'd0;
	mem_6[12] = 64'd0;
	mem_6[13] = 64'd0;
	mem_6[14] = 64'd0;
	mem_6[15] = 64'd0;
	mem_6[16] = 64'd0;
	mem_6[17] = 64'd0;
	mem_6[18] = 64'd0;
	mem_6[19] = 64'd0;
	mem_6[20] = 64'd0;
	mem_6[21] = 64'd0;
	mem_6[22] = 64'd0;
	mem_6[23] = 64'd0;
	mem_6[24] = 64'd0;
	mem_6[25] = 64'd0;
	mem_6[26] = 64'd0;
	mem_6[27] = 64'd0;
	mem_6[28] = 64'd0;
	mem_6[29] = 64'd0;
	mem_6[30] = 64'd0;
	mem_6[31] = 64'd0;
	mem_6[32] = 64'd0;
	mem_6[33] = 64'd0;
	mem_6[34] = 64'd0;
	mem_6[35] = 64'd0;
	mem_6[36] = 64'd0;
	mem_6[37] = 64'd0;
	mem_6[38] = 64'd0;
	mem_6[39] = 64'd0;
	mem_6[40] = 64'd0;
	mem_6[41] = 64'd0;
	mem_6[42] = 64'd0;
	mem_6[43] = 64'd0;
	mem_6[44] = 64'd0;
	mem_6[45] = 64'd0;
	mem_6[46] = 64'd0;
	mem_6[47] = 64'd0;
	mem_6[48] = 64'd0;
	mem_6[49] = 64'd0;
	mem_6[50] = 64'd0;
	mem_6[51] = 64'd0;
	mem_6[52] = 64'd0;
	mem_6[53] = 64'd0;
	mem_6[54] = 64'd0;
	mem_6[55] = 64'd0;
	mem_6[56] = 64'd0;
	mem_6[57] = 64'd0;
	mem_6[58] = 64'd0;
	mem_6[59] = 64'd0;
	mem_6[60] = 64'd0;
	mem_6[61] = 64'd0;
	mem_6[62] = 64'd0;
	mem_6[63] = 64'd0;
	mem_6[64] = 64'd0;
	mem_6[65] = 64'd0;
	mem_6[66] = 64'd0;
	mem_6[67] = 64'd0;
	mem_6[68] = 64'd0;
	mem_6[69] = 64'd0;
	mem_6[70] = 64'd0;
	mem_6[71] = 64'd0;
	mem_6[72] = 64'd0;
	mem_6[73] = 64'd0;
	mem_6[74] = 64'd0;
	mem_6[75] = 64'd0;
	mem_6[76] = 64'd0;
	mem_6[77] = 64'd0;
	mem_6[78] = 64'd0;
	mem_6[79] = 64'd0;
	mem_6[80] = 64'd0;
	mem_6[81] = 64'd0;
	mem_6[82] = 64'd0;
	mem_6[83] = 64'd0;
	mem_6[84] = 64'd0;
	mem_6[85] = 64'd0;
	mem_6[86] = 64'd0;
	mem_6[87] = 64'd0;
	mem_6[88] = 64'd0;
	mem_6[89] = 64'd0;
	mem_6[90] = 64'd0;
	mem_6[91] = 64'd0;
	mem_6[92] = 64'd0;
	mem_6[93] = 64'd0;
	mem_6[94] = 64'd0;
	mem_6[95] = 64'd0;
	mem_6[96] = 64'd0;
	mem_6[97] = 64'd0;
	mem_6[98] = 64'd0;
	mem_6[99] = 64'd0;
	mem_6[100] = 64'd0;
	mem_6[101] = 64'd0;
	mem_6[102] = 64'd0;
	mem_6[103] = 64'd0;
	mem_6[104] = 64'd0;
	mem_6[105] = 64'd0;
	mem_6[106] = 64'd0;
	mem_6[107] = 64'd0;
	mem_6[108] = 64'd0;
	mem_6[109] = 64'd0;
	mem_6[110] = 64'd0;
	mem_6[111] = 64'd0;
	mem_6[112] = 64'd0;
	mem_6[113] = 64'd0;
	mem_6[114] = 64'd0;
	mem_6[115] = 64'd0;
	mem_6[116] = 64'd0;
	mem_6[117] = 64'd0;
	mem_6[118] = 64'd0;
	mem_6[119] = 64'd0;
	mem_6[120] = 64'd0;
	mem_6[121] = 64'd0;
	mem_6[122] = 64'd0;
	mem_6[123] = 64'd0;
	mem_6[124] = 64'd0;
	mem_6[125] = 64'd0;
	mem_6[126] = 64'd0;
	mem_6[127] = 64'd0;
	mem_6[128] = 64'd0;
	mem_6[129] = 64'd0;
	mem_6[130] = 64'd0;
	mem_6[131] = 64'd0;
	mem_6[132] = 64'd0;
	mem_6[133] = 64'd0;
	mem_6[134] = 64'd0;
	mem_6[135] = 64'd0;
	mem_6[136] = 64'd0;
	mem_6[137] = 64'd0;
	mem_6[138] = 64'd0;
	mem_6[139] = 64'd0;
	mem_6[140] = 64'd0;
	mem_6[141] = 64'd0;
	mem_6[142] = 64'd0;
	mem_6[143] = 64'd0;
	mem_6[144] = 64'd0;
	mem_6[145] = 64'd0;
	mem_6[146] = 64'd0;
	mem_6[147] = 64'd0;
	mem_6[148] = 64'd0;
	mem_6[149] = 64'd0;
	mem_6[150] = 64'd0;
	mem_6[151] = 64'd0;
	mem_6[152] = 64'd0;
	mem_6[153] = 64'd0;
	mem_6[154] = 64'd0;
	mem_6[155] = 64'd0;
	mem_6[156] = 64'd0;
	mem_6[157] = 64'd0;
	mem_6[158] = 64'd0;
	mem_6[159] = 64'd0;
	mem_6[160] = 64'd0;
	mem_6[161] = 64'd0;
	mem_6[162] = 64'd0;
	mem_6[163] = 64'd0;
	mem_6[164] = 64'd0;
	mem_6[165] = 64'd0;
	mem_6[166] = 64'd0;
	mem_6[167] = 64'd0;
	mem_6[168] = 64'd0;
	mem_6[169] = 64'd0;
	mem_6[170] = 64'd0;
	mem_6[171] = 64'd0;
	mem_6[172] = 64'd0;
	mem_6[173] = 64'd0;
	mem_6[174] = 64'd0;
	mem_6[175] = 64'd0;
	mem_6[176] = 64'd0;
	mem_6[177] = 64'd0;
	mem_6[178] = 64'd0;
	mem_6[179] = 64'd0;
	mem_6[180] = 64'd0;
	mem_6[181] = 64'd0;
	mem_6[182] = 64'd0;
	mem_6[183] = 64'd0;
	mem_6[184] = 64'd0;
	mem_6[185] = 64'd0;
	mem_6[186] = 64'd0;
	mem_6[187] = 64'd0;
	mem_6[188] = 64'd0;
	mem_6[189] = 64'd0;
	mem_6[190] = 64'd0;
	mem_6[191] = 64'd0;
	mem_6[192] = 64'd0;
	mem_6[193] = 64'd0;
	mem_6[194] = 64'd0;
	mem_6[195] = 64'd0;
	mem_6[196] = 64'd0;
	mem_6[197] = 64'd0;
	mem_6[198] = 64'd0;
	mem_6[199] = 64'd0;
	mem_6[200] = 64'd0;
	mem_6[201] = 64'd0;
	mem_6[202] = 64'd0;
	mem_6[203] = 64'd0;
	mem_6[204] = 64'd0;
	mem_6[205] = 64'd0;
	mem_6[206] = 64'd0;
	mem_6[207] = 64'd0;
	mem_6[208] = 64'd0;
	mem_6[209] = 64'd0;
	mem_6[210] = 64'd0;
	mem_6[211] = 64'd0;
	mem_6[212] = 64'd0;
	mem_6[213] = 64'd0;
	mem_6[214] = 64'd0;
	mem_6[215] = 64'd0;
	mem_6[216] = 64'd0;
	mem_6[217] = 64'd0;
	mem_6[218] = 64'd0;
	mem_6[219] = 64'd0;
	mem_6[220] = 64'd0;
	mem_6[221] = 64'd0;
	mem_6[222] = 64'd0;
	mem_6[223] = 64'd0;
	mem_6[224] = 64'd0;
	mem_6[225] = 64'd0;
	mem_6[226] = 64'd0;
	mem_6[227] = 64'd0;
	mem_6[228] = 64'd0;
	mem_6[229] = 64'd0;
	mem_6[230] = 64'd0;
	mem_6[231] = 64'd0;
	mem_6[232] = 64'd0;
	mem_6[233] = 64'd0;
	mem_6[234] = 64'd0;
	mem_6[235] = 64'd0;
	mem_6[236] = 64'd0;
	mem_6[237] = 64'd0;
	mem_6[238] = 64'd0;
	mem_6[239] = 64'd0;
	mem_6[240] = 64'd0;
	mem_6[241] = 64'd0;
	mem_6[242] = 64'd0;
	mem_6[243] = 64'd0;
	mem_6[244] = 64'd0;
	mem_6[245] = 64'd0;
	mem_6[246] = 64'd0;
	mem_6[247] = 64'd0;
	mem_6[248] = 64'd0;
	mem_6[249] = 64'd0;
	mem_6[250] = 64'd0;
	mem_6[251] = 64'd0;
	mem_6[252] = 64'd0;
	mem_6[253] = 64'd0;
	mem_6[254] = 64'd0;
	mem_6[255] = 64'd0;
	mem_6[256] = 64'd0;
	mem_6[257] = 64'd0;
	mem_6[258] = 64'd0;
	mem_6[259] = 64'd0;
	mem_6[260] = 64'd0;
	mem_6[261] = 64'd0;
	mem_6[262] = 64'd0;
	mem_6[263] = 64'd0;
	mem_6[264] = 64'd0;
	mem_6[265] = 64'd0;
	mem_6[266] = 64'd0;
	mem_6[267] = 64'd0;
	mem_6[268] = 64'd0;
	mem_6[269] = 64'd0;
	mem_6[270] = 64'd0;
	mem_6[271] = 64'd0;
	mem_6[272] = 64'd0;
	mem_6[273] = 64'd0;
	mem_6[274] = 64'd0;
	mem_6[275] = 64'd0;
	mem_6[276] = 64'd0;
	mem_6[277] = 64'd0;
	mem_6[278] = 64'd0;
	mem_6[279] = 64'd0;
	mem_6[280] = 64'd0;
	mem_6[281] = 64'd0;
	mem_6[282] = 64'd0;
	mem_6[283] = 64'd0;
	mem_6[284] = 64'd0;
	mem_6[285] = 64'd0;
	mem_6[286] = 64'd0;
	mem_6[287] = 64'd0;
	mem_6[288] = 64'd0;
	mem_6[289] = 64'd0;
	mem_6[290] = 64'd0;
	mem_6[291] = 64'd0;
	mem_6[292] = 64'd0;
	mem_6[293] = 64'd0;
	mem_6[294] = 64'd0;
	mem_6[295] = 64'd0;
	mem_6[296] = 64'd0;
	mem_6[297] = 64'd0;
	mem_6[298] = 64'd0;
	mem_6[299] = 64'd0;
	mem_6[300] = 64'd0;
	mem_6[301] = 64'd0;
	mem_6[302] = 64'd0;
	mem_6[303] = 64'd0;
	mem_6[304] = 64'd0;
	mem_6[305] = 64'd0;
	mem_6[306] = 64'd0;
	mem_6[307] = 64'd0;
	mem_6[308] = 64'd0;
	mem_6[309] = 64'd0;
	mem_6[310] = 64'd0;
	mem_6[311] = 64'd0;
	mem_6[312] = 64'd0;
	mem_6[313] = 64'd0;
	mem_6[314] = 64'd0;
	mem_6[315] = 64'd0;
	mem_6[316] = 64'd0;
	mem_6[317] = 64'd0;
	mem_6[318] = 64'd0;
	mem_6[319] = 64'd0;
	mem_6[320] = 64'd0;
	mem_6[321] = 64'd0;
	mem_6[322] = 64'd0;
	mem_6[323] = 64'd0;
	mem_6[324] = 64'd0;
	mem_6[325] = 64'd0;
	mem_6[326] = 64'd0;
	mem_6[327] = 64'd0;
	mem_6[328] = 64'd0;
	mem_6[329] = 64'd0;
	mem_6[330] = 64'd0;
	mem_6[331] = 64'd0;
	mem_6[332] = 64'd0;
	mem_6[333] = 64'd0;
	mem_6[334] = 64'd0;
	mem_6[335] = 64'd0;
	mem_6[336] = 64'd0;
	mem_6[337] = 64'd0;
	mem_6[338] = 64'd0;
	mem_6[339] = 64'd0;
	mem_6[340] = 64'd0;
	mem_6[341] = 64'd0;
	mem_6[342] = 64'd0;
	mem_6[343] = 64'd0;
	mem_6[344] = 64'd0;
	mem_6[345] = 64'd0;
	mem_6[346] = 64'd0;
	mem_6[347] = 64'd0;
	mem_6[348] = 64'd0;
	mem_6[349] = 64'd0;
	mem_6[350] = 64'd0;
	mem_6[351] = 64'd0;
	mem_6[352] = 64'd0;
	mem_6[353] = 64'd0;
	mem_6[354] = 64'd0;
	mem_6[355] = 64'd0;
	mem_6[356] = 64'd0;
	mem_6[357] = 64'd0;
	mem_6[358] = 64'd0;
	mem_6[359] = 64'd0;
	mem_6[360] = 64'd0;
	mem_6[361] = 64'd0;
	mem_6[362] = 64'd0;
	mem_6[363] = 64'd0;
	mem_6[364] = 64'd0;
	mem_6[365] = 64'd0;
	mem_6[366] = 64'd0;
	mem_6[367] = 64'd0;
	mem_6[368] = 64'd0;
	mem_6[369] = 64'd0;
	mem_6[370] = 64'd0;
	mem_6[371] = 64'd0;
	mem_6[372] = 64'd0;
	mem_6[373] = 64'd0;
	mem_6[374] = 64'd0;
	mem_6[375] = 64'd0;
	mem_6[376] = 64'd0;
	mem_6[377] = 64'd0;
	mem_6[378] = 64'd0;
	mem_6[379] = 64'd0;
	mem_6[380] = 64'd0;
	mem_6[381] = 64'd0;
	mem_6[382] = 64'd0;
	mem_6[383] = 64'd0;
	mem_6[384] = 64'd0;
	mem_6[385] = 64'd0;
	mem_6[386] = 64'd0;
	mem_6[387] = 64'd0;
	mem_6[388] = 64'd0;
	mem_6[389] = 64'd0;
	mem_6[390] = 64'd0;
	mem_6[391] = 64'd0;
	mem_6[392] = 64'd0;
	mem_6[393] = 64'd0;
	mem_6[394] = 64'd0;
	mem_6[395] = 64'd0;
	mem_6[396] = 64'd0;
	mem_6[397] = 64'd0;
	mem_6[398] = 64'd0;
	mem_6[399] = 64'd0;
	mem_6[400] = 64'd0;
	mem_6[401] = 64'd0;
	mem_6[402] = 64'd0;
	mem_6[403] = 64'd0;
	mem_6[404] = 64'd0;
	mem_6[405] = 64'd0;
	mem_6[406] = 64'd0;
	mem_6[407] = 64'd0;
	mem_6[408] = 64'd0;
	mem_6[409] = 64'd0;
	mem_6[410] = 64'd0;
	mem_6[411] = 64'd0;
	mem_6[412] = 64'd0;
	mem_6[413] = 64'd0;
	mem_6[414] = 64'd0;
	mem_6[415] = 64'd0;
	mem_6[416] = 64'd0;
	mem_6[417] = 64'd0;
	mem_6[418] = 64'd0;
	mem_6[419] = 64'd0;
	mem_6[420] = 64'd0;
	mem_6[421] = 64'd0;
	mem_6[422] = 64'd0;
	mem_6[423] = 64'd0;
	mem_6[424] = 64'd0;
	mem_6[425] = 64'd0;
	mem_6[426] = 64'd0;
	mem_6[427] = 64'd0;
	mem_6[428] = 64'd0;
	mem_6[429] = 64'd0;
	mem_6[430] = 64'd0;
	mem_6[431] = 64'd0;
	mem_6[432] = 64'd0;
	mem_6[433] = 64'd0;
	mem_6[434] = 64'd0;
	mem_6[435] = 64'd0;
	mem_6[436] = 64'd0;
	mem_6[437] = 64'd0;
	mem_6[438] = 64'd0;
	mem_6[439] = 64'd0;
	mem_6[440] = 64'd0;
	mem_6[441] = 64'd0;
	mem_6[442] = 64'd0;
	mem_6[443] = 64'd0;
	mem_6[444] = 64'd0;
	mem_6[445] = 64'd0;
	mem_6[446] = 64'd0;
	mem_6[447] = 64'd0;
	mem_6[448] = 64'd0;
	mem_6[449] = 64'd0;
	mem_6[450] = 64'd0;
	mem_6[451] = 64'd0;
	mem_6[452] = 64'd0;
	mem_6[453] = 64'd0;
	mem_6[454] = 64'd0;
	mem_6[455] = 64'd0;
	mem_6[456] = 64'd0;
	mem_6[457] = 64'd0;
	mem_6[458] = 64'd0;
	mem_6[459] = 64'd0;
	mem_6[460] = 64'd0;
	mem_6[461] = 64'd0;
	mem_6[462] = 64'd0;
	mem_6[463] = 64'd0;
	mem_6[464] = 64'd0;
	mem_6[465] = 64'd0;
	mem_6[466] = 64'd0;
	mem_6[467] = 64'd0;
	mem_6[468] = 64'd0;
	mem_6[469] = 64'd0;
	mem_6[470] = 64'd0;
	mem_6[471] = 64'd0;
	mem_6[472] = 64'd0;
	mem_6[473] = 64'd0;
	mem_6[474] = 64'd0;
	mem_6[475] = 64'd0;
	mem_6[476] = 64'd0;
	mem_6[477] = 64'd0;
	mem_6[478] = 64'd0;
	mem_6[479] = 64'd0;
	mem_6[480] = 64'd0;
	mem_6[481] = 64'd0;
	mem_6[482] = 64'd0;
	mem_6[483] = 64'd0;
	mem_6[484] = 64'd0;
	mem_6[485] = 64'd0;
	mem_6[486] = 64'd0;
	mem_6[487] = 64'd0;
	mem_6[488] = 64'd0;
	mem_6[489] = 64'd0;
	mem_6[490] = 64'd0;
	mem_6[491] = 64'd0;
	mem_6[492] = 64'd0;
	mem_6[493] = 64'd0;
	mem_6[494] = 64'd0;
	mem_6[495] = 64'd0;
	mem_6[496] = 64'd0;
	mem_6[497] = 64'd0;
	mem_6[498] = 64'd0;
	mem_6[499] = 64'd0;
	mem_6[500] = 64'd0;
	mem_6[501] = 64'd0;
	mem_6[502] = 64'd0;
	mem_6[503] = 64'd0;
	mem_6[504] = 64'd0;
	mem_6[505] = 64'd0;
	mem_6[506] = 64'd0;
	mem_6[507] = 64'd0;
	mem_6[508] = 64'd0;
	mem_6[509] = 64'd0;
	mem_6[510] = 64'd0;
	mem_6[511] = 64'd0;
	mem_6[512] = 64'd0;
	mem_6[513] = 64'd0;
	mem_6[514] = 64'd0;
	mem_6[515] = 64'd0;
	mem_6[516] = 64'd0;
	mem_6[517] = 64'd0;
	mem_6[518] = 64'd0;
	mem_6[519] = 64'd0;
	mem_6[520] = 64'd0;
	mem_6[521] = 64'd0;
	mem_6[522] = 64'd0;
	mem_6[523] = 64'd0;
	mem_6[524] = 64'd0;
	mem_6[525] = 64'd0;
	mem_6[526] = 64'd0;
	mem_6[527] = 64'd0;
	mem_6[528] = 64'd0;
	mem_6[529] = 64'd0;
	mem_6[530] = 64'd0;
	mem_6[531] = 64'd0;
	mem_6[532] = 64'd0;
	mem_6[533] = 64'd0;
	mem_6[534] = 64'd0;
	mem_6[535] = 64'd0;
	mem_6[536] = 64'd0;
	mem_6[537] = 64'd0;
	mem_6[538] = 64'd0;
	mem_6[539] = 64'd0;
	mem_6[540] = 64'd0;
	mem_6[541] = 64'd0;
	mem_6[542] = 64'd0;
	mem_6[543] = 64'd0;
	mem_6[544] = 64'd0;
	mem_6[545] = 64'd0;
	mem_6[546] = 64'd0;
	mem_6[547] = 64'd0;
	mem_6[548] = 64'd0;
	mem_6[549] = 64'd0;
	mem_6[550] = 64'd0;
	mem_6[551] = 64'd0;
	mem_6[552] = 64'd0;
	mem_6[553] = 64'd0;
	mem_6[554] = 64'd0;
	mem_6[555] = 64'd0;
	mem_6[556] = 64'd0;
	mem_6[557] = 64'd0;
	mem_6[558] = 64'd0;
	mem_6[559] = 64'd0;
	mem_6[560] = 64'd0;
	mem_6[561] = 64'd0;
	mem_6[562] = 64'd0;
	mem_6[563] = 64'd0;
	mem_6[564] = 64'd0;
	mem_6[565] = 64'd0;
	mem_6[566] = 64'd0;
	mem_6[567] = 64'd0;
	mem_6[568] = 64'd0;
	mem_6[569] = 64'd0;
	mem_6[570] = 64'd0;
	mem_6[571] = 64'd0;
	mem_6[572] = 64'd0;
	mem_6[573] = 64'd0;
	mem_6[574] = 64'd0;
	mem_6[575] = 64'd0;
	mem_6[576] = 64'd0;
	mem_6[577] = 64'd0;
	mem_6[578] = 64'd0;
	mem_6[579] = 64'd0;
	mem_6[580] = 64'd0;
	mem_6[581] = 64'd0;
	mem_6[582] = 64'd0;
	mem_6[583] = 64'd0;
	mem_6[584] = 64'd0;
	mem_6[585] = 64'd0;
	mem_6[586] = 64'd0;
	mem_6[587] = 64'd0;
	mem_6[588] = 64'd0;
	mem_6[589] = 64'd0;
	mem_6[590] = 64'd0;
	mem_6[591] = 64'd0;
	mem_6[592] = 64'd0;
	mem_6[593] = 64'd0;
	mem_6[594] = 64'd0;
	mem_6[595] = 64'd0;
	mem_6[596] = 64'd0;
	mem_6[597] = 64'd0;
	mem_6[598] = 64'd0;
	mem_6[599] = 64'd0;
	mem_6[600] = 64'd0;
	mem_6[601] = 64'd0;
	mem_6[602] = 64'd0;
	mem_6[603] = 64'd0;
	mem_6[604] = 64'd0;
	mem_6[605] = 64'd0;
	mem_6[606] = 64'd0;
	mem_6[607] = 64'd0;
	mem_6[608] = 64'd0;
	mem_6[609] = 64'd0;
	mem_6[610] = 64'd0;
	mem_6[611] = 64'd0;
	mem_6[612] = 64'd0;
	mem_6[613] = 64'd0;
	mem_6[614] = 64'd0;
	mem_6[615] = 64'd0;
	mem_6[616] = 64'd0;
	mem_6[617] = 64'd0;
	mem_6[618] = 64'd0;
	mem_6[619] = 64'd0;
	mem_6[620] = 64'd0;
	mem_6[621] = 64'd0;
	mem_6[622] = 64'd0;
	mem_6[623] = 64'd0;
	mem_6[624] = 64'd0;
	mem_6[625] = 64'd0;
	mem_6[626] = 64'd0;
	mem_6[627] = 64'd0;
	mem_6[628] = 64'd0;
	mem_6[629] = 64'd0;
	mem_6[630] = 64'd0;
	mem_6[631] = 64'd0;
	mem_6[632] = 64'd0;
	mem_6[633] = 64'd0;
	mem_6[634] = 64'd0;
	mem_6[635] = 64'd0;
	mem_6[636] = 64'd0;
	mem_6[637] = 64'd0;
	mem_6[638] = 64'd0;
	mem_6[639] = 64'd0;
	mem_6[640] = 64'd0;
	mem_6[641] = 64'd0;
	mem_6[642] = 64'd0;
	mem_6[643] = 64'd0;
	mem_6[644] = 64'd0;
	mem_6[645] = 64'd0;
	mem_6[646] = 64'd0;
	mem_6[647] = 64'd0;
	mem_6[648] = 64'd0;
	mem_6[649] = 64'd0;
	mem_6[650] = 64'd0;
	mem_6[651] = 64'd0;
	mem_6[652] = 64'd0;
	mem_6[653] = 64'd0;
	mem_6[654] = 64'd0;
	mem_6[655] = 64'd0;
	mem_6[656] = 64'd0;
	mem_6[657] = 64'd0;
	mem_6[658] = 64'd0;
	mem_6[659] = 64'd0;
	mem_6[660] = 64'd0;
	mem_6[661] = 64'd0;
	mem_6[662] = 64'd0;
	mem_6[663] = 64'd0;
	mem_6[664] = 64'd0;
	mem_6[665] = 64'd0;
	mem_6[666] = 64'd0;
	mem_6[667] = 64'd0;
	mem_6[668] = 64'd0;
	mem_6[669] = 64'd0;
	mem_6[670] = 64'd0;
	mem_6[671] = 64'd0;
	mem_6[672] = 64'd0;
	mem_6[673] = 64'd0;
	mem_6[674] = 64'd0;
	mem_6[675] = 64'd0;
	mem_6[676] = 64'd0;
	mem_6[677] = 64'd0;
	mem_6[678] = 64'd0;
	mem_6[679] = 64'd0;
	mem_6[680] = 64'd0;
	mem_6[681] = 64'd0;
	mem_6[682] = 64'd0;
	mem_6[683] = 64'd0;
	mem_6[684] = 64'd0;
	mem_6[685] = 64'd0;
	mem_6[686] = 64'd0;
	mem_6[687] = 64'd0;
	mem_6[688] = 64'd0;
	mem_6[689] = 64'd0;
	mem_6[690] = 64'd0;
	mem_6[691] = 64'd0;
	mem_6[692] = 64'd0;
	mem_6[693] = 64'd0;
	mem_6[694] = 64'd0;
	mem_6[695] = 64'd0;
	mem_6[696] = 64'd0;
	mem_6[697] = 64'd0;
	mem_6[698] = 64'd0;
	mem_6[699] = 64'd0;
	mem_6[700] = 64'd0;
	mem_6[701] = 64'd0;
	mem_6[702] = 64'd0;
	mem_6[703] = 64'd0;
	mem_6[704] = 64'd0;
	mem_6[705] = 64'd0;
	mem_6[706] = 64'd0;
	mem_6[707] = 64'd0;
	mem_6[708] = 64'd0;
	mem_6[709] = 64'd0;
	mem_6[710] = 64'd0;
	mem_6[711] = 64'd0;
	mem_6[712] = 64'd0;
	mem_6[713] = 64'd0;
	mem_6[714] = 64'd0;
	mem_6[715] = 64'd0;
	mem_6[716] = 64'd0;
	mem_6[717] = 64'd0;
	mem_6[718] = 64'd0;
	mem_6[719] = 64'd0;
	mem_6[720] = 64'd0;
	mem_6[721] = 64'd0;
	mem_6[722] = 64'd0;
	mem_6[723] = 64'd0;
	mem_6[724] = 64'd0;
	mem_6[725] = 64'd0;
	mem_6[726] = 64'd0;
	mem_6[727] = 64'd0;
	mem_6[728] = 64'd0;
	mem_6[729] = 64'd0;
	mem_6[730] = 64'd0;
	mem_6[731] = 64'd0;
	mem_6[732] = 64'd0;
	mem_6[733] = 64'd0;
	mem_6[734] = 64'd0;
	mem_6[735] = 64'd0;
	mem_6[736] = 64'd0;
	mem_6[737] = 64'd0;
	mem_6[738] = 64'd0;
	mem_6[739] = 64'd0;
	mem_6[740] = 64'd0;
	mem_6[741] = 64'd0;
	mem_6[742] = 64'd0;
	mem_6[743] = 64'd0;
	mem_6[744] = 64'd0;
	mem_6[745] = 64'd0;
	mem_6[746] = 64'd0;
	mem_6[747] = 64'd0;
	mem_6[748] = 64'd0;
	mem_6[749] = 64'd0;
	mem_6[750] = 64'd0;
	mem_6[751] = 64'd0;
	mem_6[752] = 64'd0;
	mem_6[753] = 64'd0;
	mem_6[754] = 64'd0;
	mem_6[755] = 64'd0;
	mem_6[756] = 64'd0;
	mem_6[757] = 64'd0;
	mem_6[758] = 64'd0;
	mem_6[759] = 64'd0;
	mem_6[760] = 64'd0;
	mem_6[761] = 64'd0;
	mem_6[762] = 64'd0;
	mem_6[763] = 64'd0;
	mem_6[764] = 64'd0;
	mem_6[765] = 64'd0;
	mem_6[766] = 64'd0;
	mem_6[767] = 64'd0;
	mem_6[768] = 64'd0;
	mem_6[769] = 64'd0;
	mem_6[770] = 64'd0;
	mem_6[771] = 64'd0;
	mem_6[772] = 64'd0;
	mem_6[773] = 64'd0;
	mem_6[774] = 64'd0;
	mem_6[775] = 64'd0;
	mem_6[776] = 64'd0;
	mem_6[777] = 64'd0;
	mem_6[778] = 64'd0;
	mem_6[779] = 64'd0;
	mem_6[780] = 64'd0;
	mem_6[781] = 64'd0;
	mem_6[782] = 64'd0;
	mem_6[783] = 64'd0;
	mem_6[784] = 64'd0;
	mem_6[785] = 64'd0;
	mem_6[786] = 64'd0;
	mem_6[787] = 64'd0;
	mem_6[788] = 64'd0;
	mem_6[789] = 64'd0;
	mem_6[790] = 64'd0;
	mem_6[791] = 64'd0;
	mem_6[792] = 64'd0;
	mem_6[793] = 64'd0;
	mem_6[794] = 64'd0;
	mem_6[795] = 64'd0;
	mem_6[796] = 64'd0;
	mem_6[797] = 64'd0;
	mem_6[798] = 64'd0;
	mem_6[799] = 64'd0;
	mem_6[800] = 64'd0;
	mem_6[801] = 64'd0;
	mem_6[802] = 64'd0;
	mem_6[803] = 64'd0;
	mem_6[804] = 64'd0;
	mem_6[805] = 64'd0;
	mem_6[806] = 64'd0;
	mem_6[807] = 64'd0;
	mem_6[808] = 64'd0;
	mem_6[809] = 64'd0;
	mem_6[810] = 64'd0;
	mem_6[811] = 64'd0;
	mem_6[812] = 64'd0;
	mem_6[813] = 64'd0;
	mem_6[814] = 64'd0;
	mem_6[815] = 64'd0;
	mem_6[816] = 64'd0;
	mem_6[817] = 64'd0;
	mem_6[818] = 64'd0;
	mem_6[819] = 64'd0;
	mem_6[820] = 64'd0;
	mem_6[821] = 64'd0;
	mem_6[822] = 64'd0;
	mem_6[823] = 64'd0;
	mem_6[824] = 64'd0;
	mem_6[825] = 64'd0;
	mem_6[826] = 64'd0;
	mem_6[827] = 64'd0;
	mem_6[828] = 64'd0;
	mem_6[829] = 64'd0;
	mem_6[830] = 64'd0;
	mem_6[831] = 64'd0;
	mem_6[832] = 64'd0;
	mem_6[833] = 64'd0;
	mem_6[834] = 64'd0;
	mem_6[835] = 64'd0;
	mem_6[836] = 64'd0;
	mem_6[837] = 64'd0;
	mem_6[838] = 64'd0;
	mem_6[839] = 64'd0;
	mem_6[840] = 64'd0;
	mem_6[841] = 64'd0;
	mem_6[842] = 64'd0;
	mem_6[843] = 64'd0;
	mem_6[844] = 64'd0;
	mem_6[845] = 64'd0;
	mem_6[846] = 64'd0;
	mem_6[847] = 64'd0;
	mem_6[848] = 64'd0;
	mem_6[849] = 64'd0;
	mem_6[850] = 64'd0;
	mem_6[851] = 64'd0;
	mem_6[852] = 64'd0;
	mem_6[853] = 64'd0;
	mem_6[854] = 64'd0;
	mem_6[855] = 64'd0;
	mem_6[856] = 64'd0;
	mem_6[857] = 64'd0;
	mem_6[858] = 64'd0;
	mem_6[859] = 64'd0;
	mem_6[860] = 64'd0;
	mem_6[861] = 64'd0;
	mem_6[862] = 64'd0;
	mem_6[863] = 64'd0;
	mem_6[864] = 64'd0;
	mem_6[865] = 64'd0;
	mem_6[866] = 64'd0;
	mem_6[867] = 64'd0;
	mem_6[868] = 64'd0;
	mem_6[869] = 64'd0;
	mem_6[870] = 64'd0;
	mem_6[871] = 64'd0;
	mem_6[872] = 64'd0;
	mem_6[873] = 64'd0;
	mem_6[874] = 64'd0;
	mem_6[875] = 64'd0;
	mem_6[876] = 64'd0;
	mem_6[877] = 64'd0;
	mem_6[878] = 64'd0;
	mem_6[879] = 64'd0;
	mem_6[880] = 64'd0;
	mem_6[881] = 64'd0;
	mem_6[882] = 64'd0;
	mem_6[883] = 64'd0;
	mem_6[884] = 64'd0;
	mem_6[885] = 64'd0;
	mem_6[886] = 64'd0;
	mem_6[887] = 64'd0;
	mem_6[888] = 64'd0;
	mem_6[889] = 64'd0;
	mem_6[890] = 64'd0;
	mem_6[891] = 64'd0;
	mem_6[892] = 64'd0;
	mem_6[893] = 64'd0;
	mem_6[894] = 64'd0;
	mem_6[895] = 64'd0;
	mem_6[896] = 64'd0;
	mem_6[897] = 64'd0;
	mem_6[898] = 64'd0;
	mem_6[899] = 64'd0;
	mem_6[900] = 64'd0;
	mem_6[901] = 64'd0;
	mem_6[902] = 64'd0;
	mem_6[903] = 64'd0;
	mem_6[904] = 64'd0;
	mem_6[905] = 64'd0;
	mem_6[906] = 64'd0;
	mem_6[907] = 64'd0;
	mem_6[908] = 64'd0;
	mem_6[909] = 64'd0;
	mem_6[910] = 64'd0;
	mem_6[911] = 64'd0;
	mem_6[912] = 64'd0;
	mem_6[913] = 64'd0;
	mem_6[914] = 64'd0;
	mem_6[915] = 64'd0;
	mem_6[916] = 64'd0;
	mem_6[917] = 64'd0;
	mem_6[918] = 64'd0;
	mem_6[919] = 64'd0;
	mem_6[920] = 64'd0;
	mem_6[921] = 64'd0;
	mem_6[922] = 64'd0;
	mem_6[923] = 64'd0;
	mem_6[924] = 64'd0;
	mem_6[925] = 64'd0;
	mem_6[926] = 64'd0;
	mem_6[927] = 64'd0;
	mem_6[928] = 64'd0;
	mem_6[929] = 64'd0;
	mem_6[930] = 64'd0;
	mem_6[931] = 64'd0;
	mem_6[932] = 64'd0;
	mem_6[933] = 64'd0;
	mem_6[934] = 64'd0;
	mem_6[935] = 64'd0;
	mem_6[936] = 64'd0;
	mem_6[937] = 64'd0;
	mem_6[938] = 64'd0;
	mem_6[939] = 64'd0;
	mem_6[940] = 64'd0;
	mem_6[941] = 64'd0;
	mem_6[942] = 64'd0;
	mem_6[943] = 64'd0;
	mem_6[944] = 64'd0;
	mem_6[945] = 64'd0;
	mem_6[946] = 64'd0;
	mem_6[947] = 64'd0;
	mem_6[948] = 64'd0;
	mem_6[949] = 64'd0;
	mem_6[950] = 64'd0;
	mem_6[951] = 64'd0;
	mem_6[952] = 64'd0;
	mem_6[953] = 64'd0;
	mem_6[954] = 64'd0;
	mem_6[955] = 64'd0;
	mem_6[956] = 64'd0;
	mem_6[957] = 64'd0;
	mem_6[958] = 64'd0;
	mem_6[959] = 64'd0;
	mem_6[960] = 64'd0;
	mem_6[961] = 64'd0;
	mem_6[962] = 64'd0;
	mem_6[963] = 64'd0;
	mem_6[964] = 64'd0;
	mem_6[965] = 64'd0;
	mem_6[966] = 64'd0;
	mem_6[967] = 64'd0;
	mem_6[968] = 64'd0;
	mem_6[969] = 64'd0;
	mem_6[970] = 64'd0;
	mem_6[971] = 64'd0;
	mem_6[972] = 64'd0;
	mem_6[973] = 64'd0;
	mem_6[974] = 64'd0;
	mem_6[975] = 64'd0;
	mem_6[976] = 64'd0;
	mem_6[977] = 64'd0;
	mem_6[978] = 64'd0;
	mem_6[979] = 64'd0;
	mem_6[980] = 64'd0;
	mem_6[981] = 64'd0;
	mem_6[982] = 64'd0;
	mem_6[983] = 64'd0;
	mem_6[984] = 64'd0;
	mem_6[985] = 64'd0;
	mem_6[986] = 64'd0;
	mem_6[987] = 64'd0;
	mem_6[988] = 64'd0;
	mem_6[989] = 64'd0;
	mem_6[990] = 64'd0;
	mem_6[991] = 64'd0;
	mem_6[992] = 64'd0;
	mem_6[993] = 64'd0;
	mem_6[994] = 64'd0;
	mem_6[995] = 64'd0;
	mem_6[996] = 64'd0;
	mem_6[997] = 64'd0;
	mem_6[998] = 64'd0;
	mem_6[999] = 64'd0;
	mem_6[1000] = 64'd0;
	mem_6[1001] = 64'd0;
	mem_6[1002] = 64'd0;
	mem_6[1003] = 64'd0;
	mem_6[1004] = 64'd0;
	mem_6[1005] = 64'd0;
	mem_6[1006] = 64'd0;
	mem_6[1007] = 64'd0;
	mem_6[1008] = 64'd0;
	mem_6[1009] = 64'd0;
	mem_6[1010] = 64'd0;
	mem_6[1011] = 64'd0;
	mem_6[1012] = 64'd0;
	mem_6[1013] = 64'd0;
	mem_6[1014] = 64'd0;
	mem_6[1015] = 64'd0;
	mem_6[1016] = 64'd0;
	mem_6[1017] = 64'd0;
	mem_6[1018] = 64'd0;
	mem_6[1019] = 64'd0;
	mem_6[1020] = 64'd0;
	mem_6[1021] = 64'd0;
	mem_6[1022] = 64'd0;
	mem_6[1023] = 64'd0;
	mem_7[0] = 64'd0;
	mem_7[1] = 64'd0;
	mem_7[2] = 64'd0;
	mem_7[3] = 64'd0;
	mem_7[4] = 64'd0;
	mem_7[5] = 64'd0;
	mem_7[6] = 64'd0;
	mem_7[7] = 64'd0;
	mem_7[8] = 64'd0;
	mem_7[9] = 64'd0;
	mem_7[10] = 64'd0;
	mem_7[11] = 64'd0;
	mem_7[12] = 64'd0;
	mem_7[13] = 64'd0;
	mem_7[14] = 64'd0;
	mem_7[15] = 64'd0;
	mem_7[16] = 64'd0;
	mem_7[17] = 64'd0;
	mem_7[18] = 64'd0;
	mem_7[19] = 64'd0;
	mem_7[20] = 64'd0;
	mem_7[21] = 64'd0;
	mem_7[22] = 64'd0;
	mem_7[23] = 64'd0;
	mem_7[24] = 64'd0;
	mem_7[25] = 64'd0;
	mem_7[26] = 64'd0;
	mem_7[27] = 64'd0;
	mem_7[28] = 64'd0;
	mem_7[29] = 64'd0;
	mem_7[30] = 64'd0;
	mem_7[31] = 64'd0;
	mem_7[32] = 64'd0;
	mem_7[33] = 64'd0;
	mem_7[34] = 64'd0;
	mem_7[35] = 64'd0;
	mem_7[36] = 64'd0;
	mem_7[37] = 64'd0;
	mem_7[38] = 64'd0;
	mem_7[39] = 64'd0;
	mem_7[40] = 64'd0;
	mem_7[41] = 64'd0;
	mem_7[42] = 64'd0;
	mem_7[43] = 64'd0;
	mem_7[44] = 64'd0;
	mem_7[45] = 64'd0;
	mem_7[46] = 64'd0;
	mem_7[47] = 64'd0;
	mem_7[48] = 64'd0;
	mem_7[49] = 64'd0;
	mem_7[50] = 64'd0;
	mem_7[51] = 64'd0;
	mem_7[52] = 64'd0;
	mem_7[53] = 64'd0;
	mem_7[54] = 64'd0;
	mem_7[55] = 64'd0;
	mem_7[56] = 64'd0;
	mem_7[57] = 64'd0;
	mem_7[58] = 64'd0;
	mem_7[59] = 64'd0;
	mem_7[60] = 64'd0;
	mem_7[61] = 64'd0;
	mem_7[62] = 64'd0;
	mem_7[63] = 64'd0;
	mem_7[64] = 64'd0;
	mem_7[65] = 64'd0;
	mem_7[66] = 64'd0;
	mem_7[67] = 64'd0;
	mem_7[68] = 64'd0;
	mem_7[69] = 64'd0;
	mem_7[70] = 64'd0;
	mem_7[71] = 64'd0;
	mem_7[72] = 64'd0;
	mem_7[73] = 64'd0;
	mem_7[74] = 64'd0;
	mem_7[75] = 64'd0;
	mem_7[76] = 64'd0;
	mem_7[77] = 64'd0;
	mem_7[78] = 64'd0;
	mem_7[79] = 64'd0;
	mem_7[80] = 64'd0;
	mem_7[81] = 64'd0;
	mem_7[82] = 64'd0;
	mem_7[83] = 64'd0;
	mem_7[84] = 64'd0;
	mem_7[85] = 64'd0;
	mem_7[86] = 64'd0;
	mem_7[87] = 64'd0;
	mem_7[88] = 64'd0;
	mem_7[89] = 64'd0;
	mem_7[90] = 64'd0;
	mem_7[91] = 64'd0;
	mem_7[92] = 64'd0;
	mem_7[93] = 64'd0;
	mem_7[94] = 64'd0;
	mem_7[95] = 64'd0;
	mem_7[96] = 64'd0;
	mem_7[97] = 64'd0;
	mem_7[98] = 64'd0;
	mem_7[99] = 64'd0;
	mem_7[100] = 64'd0;
	mem_7[101] = 64'd0;
	mem_7[102] = 64'd0;
	mem_7[103] = 64'd0;
	mem_7[104] = 64'd0;
	mem_7[105] = 64'd0;
	mem_7[106] = 64'd0;
	mem_7[107] = 64'd0;
	mem_7[108] = 64'd0;
	mem_7[109] = 64'd0;
	mem_7[110] = 64'd0;
	mem_7[111] = 64'd0;
	mem_7[112] = 64'd0;
	mem_7[113] = 64'd0;
	mem_7[114] = 64'd0;
	mem_7[115] = 64'd0;
	mem_7[116] = 64'd0;
	mem_7[117] = 64'd0;
	mem_7[118] = 64'd0;
	mem_7[119] = 64'd0;
	mem_7[120] = 64'd0;
	mem_7[121] = 64'd0;
	mem_7[122] = 64'd0;
	mem_7[123] = 64'd0;
	mem_7[124] = 64'd0;
	mem_7[125] = 64'd0;
	mem_7[126] = 64'd0;
	mem_7[127] = 64'd0;
	mem_7[128] = 64'd0;
	mem_7[129] = 64'd0;
	mem_7[130] = 64'd0;
	mem_7[131] = 64'd0;
	mem_7[132] = 64'd0;
	mem_7[133] = 64'd0;
	mem_7[134] = 64'd0;
	mem_7[135] = 64'd0;
	mem_7[136] = 64'd0;
	mem_7[137] = 64'd0;
	mem_7[138] = 64'd0;
	mem_7[139] = 64'd0;
	mem_7[140] = 64'd0;
	mem_7[141] = 64'd0;
	mem_7[142] = 64'd0;
	mem_7[143] = 64'd0;
	mem_7[144] = 64'd0;
	mem_7[145] = 64'd0;
	mem_7[146] = 64'd0;
	mem_7[147] = 64'd0;
	mem_7[148] = 64'd0;
	mem_7[149] = 64'd0;
	mem_7[150] = 64'd0;
	mem_7[151] = 64'd0;
	mem_7[152] = 64'd0;
	mem_7[153] = 64'd0;
	mem_7[154] = 64'd0;
	mem_7[155] = 64'd0;
	mem_7[156] = 64'd0;
	mem_7[157] = 64'd0;
	mem_7[158] = 64'd0;
	mem_7[159] = 64'd0;
	mem_7[160] = 64'd0;
	mem_7[161] = 64'd0;
	mem_7[162] = 64'd0;
	mem_7[163] = 64'd0;
	mem_7[164] = 64'd0;
	mem_7[165] = 64'd0;
	mem_7[166] = 64'd0;
	mem_7[167] = 64'd0;
	mem_7[168] = 64'd0;
	mem_7[169] = 64'd0;
	mem_7[170] = 64'd0;
	mem_7[171] = 64'd0;
	mem_7[172] = 64'd0;
	mem_7[173] = 64'd0;
	mem_7[174] = 64'd0;
	mem_7[175] = 64'd0;
	mem_7[176] = 64'd0;
	mem_7[177] = 64'd0;
	mem_7[178] = 64'd0;
	mem_7[179] = 64'd0;
	mem_7[180] = 64'd0;
	mem_7[181] = 64'd0;
	mem_7[182] = 64'd0;
	mem_7[183] = 64'd0;
	mem_7[184] = 64'd0;
	mem_7[185] = 64'd0;
	mem_7[186] = 64'd0;
	mem_7[187] = 64'd0;
	mem_7[188] = 64'd0;
	mem_7[189] = 64'd0;
	mem_7[190] = 64'd0;
	mem_7[191] = 64'd0;
	mem_7[192] = 64'd0;
	mem_7[193] = 64'd0;
	mem_7[194] = 64'd0;
	mem_7[195] = 64'd0;
	mem_7[196] = 64'd0;
	mem_7[197] = 64'd0;
	mem_7[198] = 64'd0;
	mem_7[199] = 64'd0;
	mem_7[200] = 64'd0;
	mem_7[201] = 64'd0;
	mem_7[202] = 64'd0;
	mem_7[203] = 64'd0;
	mem_7[204] = 64'd0;
	mem_7[205] = 64'd0;
	mem_7[206] = 64'd0;
	mem_7[207] = 64'd0;
	mem_7[208] = 64'd0;
	mem_7[209] = 64'd0;
	mem_7[210] = 64'd0;
	mem_7[211] = 64'd0;
	mem_7[212] = 64'd0;
	mem_7[213] = 64'd0;
	mem_7[214] = 64'd0;
	mem_7[215] = 64'd0;
	mem_7[216] = 64'd0;
	mem_7[217] = 64'd0;
	mem_7[218] = 64'd0;
	mem_7[219] = 64'd0;
	mem_7[220] = 64'd0;
	mem_7[221] = 64'd0;
	mem_7[222] = 64'd0;
	mem_7[223] = 64'd0;
	mem_7[224] = 64'd0;
	mem_7[225] = 64'd0;
	mem_7[226] = 64'd0;
	mem_7[227] = 64'd0;
	mem_7[228] = 64'd0;
	mem_7[229] = 64'd0;
	mem_7[230] = 64'd0;
	mem_7[231] = 64'd0;
	mem_7[232] = 64'd0;
	mem_7[233] = 64'd0;
	mem_7[234] = 64'd0;
	mem_7[235] = 64'd0;
	mem_7[236] = 64'd0;
	mem_7[237] = 64'd0;
	mem_7[238] = 64'd0;
	mem_7[239] = 64'd0;
	mem_7[240] = 64'd0;
	mem_7[241] = 64'd0;
	mem_7[242] = 64'd0;
	mem_7[243] = 64'd0;
	mem_7[244] = 64'd0;
	mem_7[245] = 64'd0;
	mem_7[246] = 64'd0;
	mem_7[247] = 64'd0;
	mem_7[248] = 64'd0;
	mem_7[249] = 64'd0;
	mem_7[250] = 64'd0;
	mem_7[251] = 64'd0;
	mem_7[252] = 64'd0;
	mem_7[253] = 64'd0;
	mem_7[254] = 64'd0;
	mem_7[255] = 64'd0;
	mem_7[256] = 64'd0;
	mem_7[257] = 64'd0;
	mem_7[258] = 64'd0;
	mem_7[259] = 64'd0;
	mem_7[260] = 64'd0;
	mem_7[261] = 64'd0;
	mem_7[262] = 64'd0;
	mem_7[263] = 64'd0;
	mem_7[264] = 64'd0;
	mem_7[265] = 64'd0;
	mem_7[266] = 64'd0;
	mem_7[267] = 64'd0;
	mem_7[268] = 64'd0;
	mem_7[269] = 64'd0;
	mem_7[270] = 64'd0;
	mem_7[271] = 64'd0;
	mem_7[272] = 64'd0;
	mem_7[273] = 64'd0;
	mem_7[274] = 64'd0;
	mem_7[275] = 64'd0;
	mem_7[276] = 64'd0;
	mem_7[277] = 64'd0;
	mem_7[278] = 64'd0;
	mem_7[279] = 64'd0;
	mem_7[280] = 64'd0;
	mem_7[281] = 64'd0;
	mem_7[282] = 64'd0;
	mem_7[283] = 64'd0;
	mem_7[284] = 64'd0;
	mem_7[285] = 64'd0;
	mem_7[286] = 64'd0;
	mem_7[287] = 64'd0;
	mem_7[288] = 64'd0;
	mem_7[289] = 64'd0;
	mem_7[290] = 64'd0;
	mem_7[291] = 64'd0;
	mem_7[292] = 64'd0;
	mem_7[293] = 64'd0;
	mem_7[294] = 64'd0;
	mem_7[295] = 64'd0;
	mem_7[296] = 64'd0;
	mem_7[297] = 64'd0;
	mem_7[298] = 64'd0;
	mem_7[299] = 64'd0;
	mem_7[300] = 64'd0;
	mem_7[301] = 64'd0;
	mem_7[302] = 64'd0;
	mem_7[303] = 64'd0;
	mem_7[304] = 64'd0;
	mem_7[305] = 64'd0;
	mem_7[306] = 64'd0;
	mem_7[307] = 64'd0;
	mem_7[308] = 64'd0;
	mem_7[309] = 64'd0;
	mem_7[310] = 64'd0;
	mem_7[311] = 64'd0;
	mem_7[312] = 64'd0;
	mem_7[313] = 64'd0;
	mem_7[314] = 64'd0;
	mem_7[315] = 64'd0;
	mem_7[316] = 64'd0;
	mem_7[317] = 64'd0;
	mem_7[318] = 64'd0;
	mem_7[319] = 64'd0;
	mem_7[320] = 64'd0;
	mem_7[321] = 64'd0;
	mem_7[322] = 64'd0;
	mem_7[323] = 64'd0;
	mem_7[324] = 64'd0;
	mem_7[325] = 64'd0;
	mem_7[326] = 64'd0;
	mem_7[327] = 64'd0;
	mem_7[328] = 64'd0;
	mem_7[329] = 64'd0;
	mem_7[330] = 64'd0;
	mem_7[331] = 64'd0;
	mem_7[332] = 64'd0;
	mem_7[333] = 64'd0;
	mem_7[334] = 64'd0;
	mem_7[335] = 64'd0;
	mem_7[336] = 64'd0;
	mem_7[337] = 64'd0;
	mem_7[338] = 64'd0;
	mem_7[339] = 64'd0;
	mem_7[340] = 64'd0;
	mem_7[341] = 64'd0;
	mem_7[342] = 64'd0;
	mem_7[343] = 64'd0;
	mem_7[344] = 64'd0;
	mem_7[345] = 64'd0;
	mem_7[346] = 64'd0;
	mem_7[347] = 64'd0;
	mem_7[348] = 64'd0;
	mem_7[349] = 64'd0;
	mem_7[350] = 64'd0;
	mem_7[351] = 64'd0;
	mem_7[352] = 64'd0;
	mem_7[353] = 64'd0;
	mem_7[354] = 64'd0;
	mem_7[355] = 64'd0;
	mem_7[356] = 64'd0;
	mem_7[357] = 64'd0;
	mem_7[358] = 64'd0;
	mem_7[359] = 64'd0;
	mem_7[360] = 64'd0;
	mem_7[361] = 64'd0;
	mem_7[362] = 64'd0;
	mem_7[363] = 64'd0;
	mem_7[364] = 64'd0;
	mem_7[365] = 64'd0;
	mem_7[366] = 64'd0;
	mem_7[367] = 64'd0;
	mem_7[368] = 64'd0;
	mem_7[369] = 64'd0;
	mem_7[370] = 64'd0;
	mem_7[371] = 64'd0;
	mem_7[372] = 64'd0;
	mem_7[373] = 64'd0;
	mem_7[374] = 64'd0;
	mem_7[375] = 64'd0;
	mem_7[376] = 64'd0;
	mem_7[377] = 64'd0;
	mem_7[378] = 64'd0;
	mem_7[379] = 64'd0;
	mem_7[380] = 64'd0;
	mem_7[381] = 64'd0;
	mem_7[382] = 64'd0;
	mem_7[383] = 64'd0;
	mem_7[384] = 64'd0;
	mem_7[385] = 64'd0;
	mem_7[386] = 64'd0;
	mem_7[387] = 64'd0;
	mem_7[388] = 64'd0;
	mem_7[389] = 64'd0;
	mem_7[390] = 64'd0;
	mem_7[391] = 64'd0;
	mem_7[392] = 64'd0;
	mem_7[393] = 64'd0;
	mem_7[394] = 64'd0;
	mem_7[395] = 64'd0;
	mem_7[396] = 64'd0;
	mem_7[397] = 64'd0;
	mem_7[398] = 64'd0;
	mem_7[399] = 64'd0;
	mem_7[400] = 64'd0;
	mem_7[401] = 64'd0;
	mem_7[402] = 64'd0;
	mem_7[403] = 64'd0;
	mem_7[404] = 64'd0;
	mem_7[405] = 64'd0;
	mem_7[406] = 64'd0;
	mem_7[407] = 64'd0;
	mem_7[408] = 64'd0;
	mem_7[409] = 64'd0;
	mem_7[410] = 64'd0;
	mem_7[411] = 64'd0;
	mem_7[412] = 64'd0;
	mem_7[413] = 64'd0;
	mem_7[414] = 64'd0;
	mem_7[415] = 64'd0;
	mem_7[416] = 64'd0;
	mem_7[417] = 64'd0;
	mem_7[418] = 64'd0;
	mem_7[419] = 64'd0;
	mem_7[420] = 64'd0;
	mem_7[421] = 64'd0;
	mem_7[422] = 64'd0;
	mem_7[423] = 64'd0;
	mem_7[424] = 64'd0;
	mem_7[425] = 64'd0;
	mem_7[426] = 64'd0;
	mem_7[427] = 64'd0;
	mem_7[428] = 64'd0;
	mem_7[429] = 64'd0;
	mem_7[430] = 64'd0;
	mem_7[431] = 64'd0;
	mem_7[432] = 64'd0;
	mem_7[433] = 64'd0;
	mem_7[434] = 64'd0;
	mem_7[435] = 64'd0;
	mem_7[436] = 64'd0;
	mem_7[437] = 64'd0;
	mem_7[438] = 64'd0;
	mem_7[439] = 64'd0;
	mem_7[440] = 64'd0;
	mem_7[441] = 64'd0;
	mem_7[442] = 64'd0;
	mem_7[443] = 64'd0;
	mem_7[444] = 64'd0;
	mem_7[445] = 64'd0;
	mem_7[446] = 64'd0;
	mem_7[447] = 64'd0;
	mem_7[448] = 64'd0;
	mem_7[449] = 64'd0;
	mem_7[450] = 64'd0;
	mem_7[451] = 64'd0;
	mem_7[452] = 64'd0;
	mem_7[453] = 64'd0;
	mem_7[454] = 64'd0;
	mem_7[455] = 64'd0;
	mem_7[456] = 64'd0;
	mem_7[457] = 64'd0;
	mem_7[458] = 64'd0;
	mem_7[459] = 64'd0;
	mem_7[460] = 64'd0;
	mem_7[461] = 64'd0;
	mem_7[462] = 64'd0;
	mem_7[463] = 64'd0;
	mem_7[464] = 64'd0;
	mem_7[465] = 64'd0;
	mem_7[466] = 64'd0;
	mem_7[467] = 64'd0;
	mem_7[468] = 64'd0;
	mem_7[469] = 64'd0;
	mem_7[470] = 64'd0;
	mem_7[471] = 64'd0;
	mem_7[472] = 64'd0;
	mem_7[473] = 64'd0;
	mem_7[474] = 64'd0;
	mem_7[475] = 64'd0;
	mem_7[476] = 64'd0;
	mem_7[477] = 64'd0;
	mem_7[478] = 64'd0;
	mem_7[479] = 64'd0;
	mem_7[480] = 64'd0;
	mem_7[481] = 64'd0;
	mem_7[482] = 64'd0;
	mem_7[483] = 64'd0;
	mem_7[484] = 64'd0;
	mem_7[485] = 64'd0;
	mem_7[486] = 64'd0;
	mem_7[487] = 64'd0;
	mem_7[488] = 64'd0;
	mem_7[489] = 64'd0;
	mem_7[490] = 64'd0;
	mem_7[491] = 64'd0;
	mem_7[492] = 64'd0;
	mem_7[493] = 64'd0;
	mem_7[494] = 64'd0;
	mem_7[495] = 64'd0;
	mem_7[496] = 64'd0;
	mem_7[497] = 64'd0;
	mem_7[498] = 64'd0;
	mem_7[499] = 64'd0;
	mem_7[500] = 64'd0;
	mem_7[501] = 64'd0;
	mem_7[502] = 64'd0;
	mem_7[503] = 64'd0;
	mem_7[504] = 64'd0;
	mem_7[505] = 64'd0;
	mem_7[506] = 64'd0;
	mem_7[507] = 64'd0;
	mem_7[508] = 64'd0;
	mem_7[509] = 64'd0;
	mem_7[510] = 64'd0;
	mem_7[511] = 64'd0;
	mem_7[512] = 64'd0;
	mem_7[513] = 64'd0;
	mem_7[514] = 64'd0;
	mem_7[515] = 64'd0;
	mem_7[516] = 64'd0;
	mem_7[517] = 64'd0;
	mem_7[518] = 64'd0;
	mem_7[519] = 64'd0;
	mem_7[520] = 64'd0;
	mem_7[521] = 64'd0;
	mem_7[522] = 64'd0;
	mem_7[523] = 64'd0;
	mem_7[524] = 64'd0;
	mem_7[525] = 64'd0;
	mem_7[526] = 64'd0;
	mem_7[527] = 64'd0;
	mem_7[528] = 64'd0;
	mem_7[529] = 64'd0;
	mem_7[530] = 64'd0;
	mem_7[531] = 64'd0;
	mem_7[532] = 64'd0;
	mem_7[533] = 64'd0;
	mem_7[534] = 64'd0;
	mem_7[535] = 64'd0;
	mem_7[536] = 64'd0;
	mem_7[537] = 64'd0;
	mem_7[538] = 64'd0;
	mem_7[539] = 64'd0;
	mem_7[540] = 64'd0;
	mem_7[541] = 64'd0;
	mem_7[542] = 64'd0;
	mem_7[543] = 64'd0;
	mem_7[544] = 64'd0;
	mem_7[545] = 64'd0;
	mem_7[546] = 64'd0;
	mem_7[547] = 64'd0;
	mem_7[548] = 64'd0;
	mem_7[549] = 64'd0;
	mem_7[550] = 64'd0;
	mem_7[551] = 64'd0;
	mem_7[552] = 64'd0;
	mem_7[553] = 64'd0;
	mem_7[554] = 64'd0;
	mem_7[555] = 64'd0;
	mem_7[556] = 64'd0;
	mem_7[557] = 64'd0;
	mem_7[558] = 64'd0;
	mem_7[559] = 64'd0;
	mem_7[560] = 64'd0;
	mem_7[561] = 64'd0;
	mem_7[562] = 64'd0;
	mem_7[563] = 64'd0;
	mem_7[564] = 64'd0;
	mem_7[565] = 64'd0;
	mem_7[566] = 64'd0;
	mem_7[567] = 64'd0;
	mem_7[568] = 64'd0;
	mem_7[569] = 64'd0;
	mem_7[570] = 64'd0;
	mem_7[571] = 64'd0;
	mem_7[572] = 64'd0;
	mem_7[573] = 64'd0;
	mem_7[574] = 64'd0;
	mem_7[575] = 64'd0;
	mem_7[576] = 64'd0;
	mem_7[577] = 64'd0;
	mem_7[578] = 64'd0;
	mem_7[579] = 64'd0;
	mem_7[580] = 64'd0;
	mem_7[581] = 64'd0;
	mem_7[582] = 64'd0;
	mem_7[583] = 64'd0;
	mem_7[584] = 64'd0;
	mem_7[585] = 64'd0;
	mem_7[586] = 64'd0;
	mem_7[587] = 64'd0;
	mem_7[588] = 64'd0;
	mem_7[589] = 64'd0;
	mem_7[590] = 64'd0;
	mem_7[591] = 64'd0;
	mem_7[592] = 64'd0;
	mem_7[593] = 64'd0;
	mem_7[594] = 64'd0;
	mem_7[595] = 64'd0;
	mem_7[596] = 64'd0;
	mem_7[597] = 64'd0;
	mem_7[598] = 64'd0;
	mem_7[599] = 64'd0;
	mem_7[600] = 64'd0;
	mem_7[601] = 64'd0;
	mem_7[602] = 64'd0;
	mem_7[603] = 64'd0;
	mem_7[604] = 64'd0;
	mem_7[605] = 64'd0;
	mem_7[606] = 64'd0;
	mem_7[607] = 64'd0;
	mem_7[608] = 64'd0;
	mem_7[609] = 64'd0;
	mem_7[610] = 64'd0;
	mem_7[611] = 64'd0;
	mem_7[612] = 64'd0;
	mem_7[613] = 64'd0;
	mem_7[614] = 64'd0;
	mem_7[615] = 64'd0;
	mem_7[616] = 64'd0;
	mem_7[617] = 64'd0;
	mem_7[618] = 64'd0;
	mem_7[619] = 64'd0;
	mem_7[620] = 64'd0;
	mem_7[621] = 64'd0;
	mem_7[622] = 64'd0;
	mem_7[623] = 64'd0;
	mem_7[624] = 64'd0;
	mem_7[625] = 64'd0;
	mem_7[626] = 64'd0;
	mem_7[627] = 64'd0;
	mem_7[628] = 64'd0;
	mem_7[629] = 64'd0;
	mem_7[630] = 64'd0;
	mem_7[631] = 64'd0;
	mem_7[632] = 64'd0;
	mem_7[633] = 64'd0;
	mem_7[634] = 64'd0;
	mem_7[635] = 64'd0;
	mem_7[636] = 64'd0;
	mem_7[637] = 64'd0;
	mem_7[638] = 64'd0;
	mem_7[639] = 64'd0;
	mem_7[640] = 64'd0;
	mem_7[641] = 64'd0;
	mem_7[642] = 64'd0;
	mem_7[643] = 64'd0;
	mem_7[644] = 64'd0;
	mem_7[645] = 64'd0;
	mem_7[646] = 64'd0;
	mem_7[647] = 64'd0;
	mem_7[648] = 64'd0;
	mem_7[649] = 64'd0;
	mem_7[650] = 64'd0;
	mem_7[651] = 64'd0;
	mem_7[652] = 64'd0;
	mem_7[653] = 64'd0;
	mem_7[654] = 64'd0;
	mem_7[655] = 64'd0;
	mem_7[656] = 64'd0;
	mem_7[657] = 64'd0;
	mem_7[658] = 64'd0;
	mem_7[659] = 64'd0;
	mem_7[660] = 64'd0;
	mem_7[661] = 64'd0;
	mem_7[662] = 64'd0;
	mem_7[663] = 64'd0;
	mem_7[664] = 64'd0;
	mem_7[665] = 64'd0;
	mem_7[666] = 64'd0;
	mem_7[667] = 64'd0;
	mem_7[668] = 64'd0;
	mem_7[669] = 64'd0;
	mem_7[670] = 64'd0;
	mem_7[671] = 64'd0;
	mem_7[672] = 64'd0;
	mem_7[673] = 64'd0;
	mem_7[674] = 64'd0;
	mem_7[675] = 64'd0;
	mem_7[676] = 64'd0;
	mem_7[677] = 64'd0;
	mem_7[678] = 64'd0;
	mem_7[679] = 64'd0;
	mem_7[680] = 64'd0;
	mem_7[681] = 64'd0;
	mem_7[682] = 64'd0;
	mem_7[683] = 64'd0;
	mem_7[684] = 64'd0;
	mem_7[685] = 64'd0;
	mem_7[686] = 64'd0;
	mem_7[687] = 64'd0;
	mem_7[688] = 64'd0;
	mem_7[689] = 64'd0;
	mem_7[690] = 64'd0;
	mem_7[691] = 64'd0;
	mem_7[692] = 64'd0;
	mem_7[693] = 64'd0;
	mem_7[694] = 64'd0;
	mem_7[695] = 64'd0;
	mem_7[696] = 64'd0;
	mem_7[697] = 64'd0;
	mem_7[698] = 64'd0;
	mem_7[699] = 64'd0;
	mem_7[700] = 64'd0;
	mem_7[701] = 64'd0;
	mem_7[702] = 64'd0;
	mem_7[703] = 64'd0;
	mem_7[704] = 64'd0;
	mem_7[705] = 64'd0;
	mem_7[706] = 64'd0;
	mem_7[707] = 64'd0;
	mem_7[708] = 64'd0;
	mem_7[709] = 64'd0;
	mem_7[710] = 64'd0;
	mem_7[711] = 64'd0;
	mem_7[712] = 64'd0;
	mem_7[713] = 64'd0;
	mem_7[714] = 64'd0;
	mem_7[715] = 64'd0;
	mem_7[716] = 64'd0;
	mem_7[717] = 64'd0;
	mem_7[718] = 64'd0;
	mem_7[719] = 64'd0;
	mem_7[720] = 64'd0;
	mem_7[721] = 64'd0;
	mem_7[722] = 64'd0;
	mem_7[723] = 64'd0;
	mem_7[724] = 64'd0;
	mem_7[725] = 64'd0;
	mem_7[726] = 64'd0;
	mem_7[727] = 64'd0;
	mem_7[728] = 64'd0;
	mem_7[729] = 64'd0;
	mem_7[730] = 64'd0;
	mem_7[731] = 64'd0;
	mem_7[732] = 64'd0;
	mem_7[733] = 64'd0;
	mem_7[734] = 64'd0;
	mem_7[735] = 64'd0;
	mem_7[736] = 64'd0;
	mem_7[737] = 64'd0;
	mem_7[738] = 64'd0;
	mem_7[739] = 64'd0;
	mem_7[740] = 64'd0;
	mem_7[741] = 64'd0;
	mem_7[742] = 64'd0;
	mem_7[743] = 64'd0;
	mem_7[744] = 64'd0;
	mem_7[745] = 64'd0;
	mem_7[746] = 64'd0;
	mem_7[747] = 64'd0;
	mem_7[748] = 64'd0;
	mem_7[749] = 64'd0;
	mem_7[750] = 64'd0;
	mem_7[751] = 64'd0;
	mem_7[752] = 64'd0;
	mem_7[753] = 64'd0;
	mem_7[754] = 64'd0;
	mem_7[755] = 64'd0;
	mem_7[756] = 64'd0;
	mem_7[757] = 64'd0;
	mem_7[758] = 64'd0;
	mem_7[759] = 64'd0;
	mem_7[760] = 64'd0;
	mem_7[761] = 64'd0;
	mem_7[762] = 64'd0;
	mem_7[763] = 64'd0;
	mem_7[764] = 64'd0;
	mem_7[765] = 64'd0;
	mem_7[766] = 64'd0;
	mem_7[767] = 64'd0;
	mem_7[768] = 64'd0;
	mem_7[769] = 64'd0;
	mem_7[770] = 64'd0;
	mem_7[771] = 64'd0;
	mem_7[772] = 64'd0;
	mem_7[773] = 64'd0;
	mem_7[774] = 64'd0;
	mem_7[775] = 64'd0;
	mem_7[776] = 64'd0;
	mem_7[777] = 64'd0;
	mem_7[778] = 64'd0;
	mem_7[779] = 64'd0;
	mem_7[780] = 64'd0;
	mem_7[781] = 64'd0;
	mem_7[782] = 64'd0;
	mem_7[783] = 64'd0;
	mem_7[784] = 64'd0;
	mem_7[785] = 64'd0;
	mem_7[786] = 64'd0;
	mem_7[787] = 64'd0;
	mem_7[788] = 64'd0;
	mem_7[789] = 64'd0;
	mem_7[790] = 64'd0;
	mem_7[791] = 64'd0;
	mem_7[792] = 64'd0;
	mem_7[793] = 64'd0;
	mem_7[794] = 64'd0;
	mem_7[795] = 64'd0;
	mem_7[796] = 64'd0;
	mem_7[797] = 64'd0;
	mem_7[798] = 64'd0;
	mem_7[799] = 64'd0;
	mem_7[800] = 64'd0;
	mem_7[801] = 64'd0;
	mem_7[802] = 64'd0;
	mem_7[803] = 64'd0;
	mem_7[804] = 64'd0;
	mem_7[805] = 64'd0;
	mem_7[806] = 64'd0;
	mem_7[807] = 64'd0;
	mem_7[808] = 64'd0;
	mem_7[809] = 64'd0;
	mem_7[810] = 64'd0;
	mem_7[811] = 64'd0;
	mem_7[812] = 64'd0;
	mem_7[813] = 64'd0;
	mem_7[814] = 64'd0;
	mem_7[815] = 64'd0;
	mem_7[816] = 64'd0;
	mem_7[817] = 64'd0;
	mem_7[818] = 64'd0;
	mem_7[819] = 64'd0;
	mem_7[820] = 64'd0;
	mem_7[821] = 64'd0;
	mem_7[822] = 64'd0;
	mem_7[823] = 64'd0;
	mem_7[824] = 64'd0;
	mem_7[825] = 64'd0;
	mem_7[826] = 64'd0;
	mem_7[827] = 64'd0;
	mem_7[828] = 64'd0;
	mem_7[829] = 64'd0;
	mem_7[830] = 64'd0;
	mem_7[831] = 64'd0;
	mem_7[832] = 64'd0;
	mem_7[833] = 64'd0;
	mem_7[834] = 64'd0;
	mem_7[835] = 64'd0;
	mem_7[836] = 64'd0;
	mem_7[837] = 64'd0;
	mem_7[838] = 64'd0;
	mem_7[839] = 64'd0;
	mem_7[840] = 64'd0;
	mem_7[841] = 64'd0;
	mem_7[842] = 64'd0;
	mem_7[843] = 64'd0;
	mem_7[844] = 64'd0;
	mem_7[845] = 64'd0;
	mem_7[846] = 64'd0;
	mem_7[847] = 64'd0;
	mem_7[848] = 64'd0;
	mem_7[849] = 64'd0;
	mem_7[850] = 64'd0;
	mem_7[851] = 64'd0;
	mem_7[852] = 64'd0;
	mem_7[853] = 64'd0;
	mem_7[854] = 64'd0;
	mem_7[855] = 64'd0;
	mem_7[856] = 64'd0;
	mem_7[857] = 64'd0;
	mem_7[858] = 64'd0;
	mem_7[859] = 64'd0;
	mem_7[860] = 64'd0;
	mem_7[861] = 64'd0;
	mem_7[862] = 64'd0;
	mem_7[863] = 64'd0;
	mem_7[864] = 64'd0;
	mem_7[865] = 64'd0;
	mem_7[866] = 64'd0;
	mem_7[867] = 64'd0;
	mem_7[868] = 64'd0;
	mem_7[869] = 64'd0;
	mem_7[870] = 64'd0;
	mem_7[871] = 64'd0;
	mem_7[872] = 64'd0;
	mem_7[873] = 64'd0;
	mem_7[874] = 64'd0;
	mem_7[875] = 64'd0;
	mem_7[876] = 64'd0;
	mem_7[877] = 64'd0;
	mem_7[878] = 64'd0;
	mem_7[879] = 64'd0;
	mem_7[880] = 64'd0;
	mem_7[881] = 64'd0;
	mem_7[882] = 64'd0;
	mem_7[883] = 64'd0;
	mem_7[884] = 64'd0;
	mem_7[885] = 64'd0;
	mem_7[886] = 64'd0;
	mem_7[887] = 64'd0;
	mem_7[888] = 64'd0;
	mem_7[889] = 64'd0;
	mem_7[890] = 64'd0;
	mem_7[891] = 64'd0;
	mem_7[892] = 64'd0;
	mem_7[893] = 64'd0;
	mem_7[894] = 64'd0;
	mem_7[895] = 64'd0;
	mem_7[896] = 64'd0;
	mem_7[897] = 64'd0;
	mem_7[898] = 64'd0;
	mem_7[899] = 64'd0;
	mem_7[900] = 64'd0;
	mem_7[901] = 64'd0;
	mem_7[902] = 64'd0;
	mem_7[903] = 64'd0;
	mem_7[904] = 64'd0;
	mem_7[905] = 64'd0;
	mem_7[906] = 64'd0;
	mem_7[907] = 64'd0;
	mem_7[908] = 64'd0;
	mem_7[909] = 64'd0;
	mem_7[910] = 64'd0;
	mem_7[911] = 64'd0;
	mem_7[912] = 64'd0;
	mem_7[913] = 64'd0;
	mem_7[914] = 64'd0;
	mem_7[915] = 64'd0;
	mem_7[916] = 64'd0;
	mem_7[917] = 64'd0;
	mem_7[918] = 64'd0;
	mem_7[919] = 64'd0;
	mem_7[920] = 64'd0;
	mem_7[921] = 64'd0;
	mem_7[922] = 64'd0;
	mem_7[923] = 64'd0;
	mem_7[924] = 64'd0;
	mem_7[925] = 64'd0;
	mem_7[926] = 64'd0;
	mem_7[927] = 64'd0;
	mem_7[928] = 64'd0;
	mem_7[929] = 64'd0;
	mem_7[930] = 64'd0;
	mem_7[931] = 64'd0;
	mem_7[932] = 64'd0;
	mem_7[933] = 64'd0;
	mem_7[934] = 64'd0;
	mem_7[935] = 64'd0;
	mem_7[936] = 64'd0;
	mem_7[937] = 64'd0;
	mem_7[938] = 64'd0;
	mem_7[939] = 64'd0;
	mem_7[940] = 64'd0;
	mem_7[941] = 64'd0;
	mem_7[942] = 64'd0;
	mem_7[943] = 64'd0;
	mem_7[944] = 64'd0;
	mem_7[945] = 64'd0;
	mem_7[946] = 64'd0;
	mem_7[947] = 64'd0;
	mem_7[948] = 64'd0;
	mem_7[949] = 64'd0;
	mem_7[950] = 64'd0;
	mem_7[951] = 64'd0;
	mem_7[952] = 64'd0;
	mem_7[953] = 64'd0;
	mem_7[954] = 64'd0;
	mem_7[955] = 64'd0;
	mem_7[956] = 64'd0;
	mem_7[957] = 64'd0;
	mem_7[958] = 64'd0;
	mem_7[959] = 64'd0;
	mem_7[960] = 64'd0;
	mem_7[961] = 64'd0;
	mem_7[962] = 64'd0;
	mem_7[963] = 64'd0;
	mem_7[964] = 64'd0;
	mem_7[965] = 64'd0;
	mem_7[966] = 64'd0;
	mem_7[967] = 64'd0;
	mem_7[968] = 64'd0;
	mem_7[969] = 64'd0;
	mem_7[970] = 64'd0;
	mem_7[971] = 64'd0;
	mem_7[972] = 64'd0;
	mem_7[973] = 64'd0;
	mem_7[974] = 64'd0;
	mem_7[975] = 64'd0;
	mem_7[976] = 64'd0;
	mem_7[977] = 64'd0;
	mem_7[978] = 64'd0;
	mem_7[979] = 64'd0;
	mem_7[980] = 64'd0;
	mem_7[981] = 64'd0;
	mem_7[982] = 64'd0;
	mem_7[983] = 64'd0;
	mem_7[984] = 64'd0;
	mem_7[985] = 64'd0;
	mem_7[986] = 64'd0;
	mem_7[987] = 64'd0;
	mem_7[988] = 64'd0;
	mem_7[989] = 64'd0;
	mem_7[990] = 64'd0;
	mem_7[991] = 64'd0;
	mem_7[992] = 64'd0;
	mem_7[993] = 64'd0;
	mem_7[994] = 64'd0;
	mem_7[995] = 64'd0;
	mem_7[996] = 64'd0;
	mem_7[997] = 64'd0;
	mem_7[998] = 64'd0;
	mem_7[999] = 64'd0;
	mem_7[1000] = 64'd0;
	mem_7[1001] = 64'd0;
	mem_7[1002] = 64'd0;
	mem_7[1003] = 64'd0;
	mem_7[1004] = 64'd0;
	mem_7[1005] = 64'd0;
	mem_7[1006] = 64'd0;
	mem_7[1007] = 64'd0;
	mem_7[1008] = 64'd0;
	mem_7[1009] = 64'd0;
	mem_7[1010] = 64'd0;
	mem_7[1011] = 64'd0;
	mem_7[1012] = 64'd0;
	mem_7[1013] = 64'd0;
	mem_7[1014] = 64'd0;
	mem_7[1015] = 64'd0;
	mem_7[1016] = 64'd0;
	mem_7[1017] = 64'd0;
	mem_7[1018] = 64'd0;
	mem_7[1019] = 64'd0;
	mem_7[1020] = 64'd0;
	mem_7[1021] = 64'd0;
	mem_7[1022] = 64'd0;
	mem_7[1023] = 64'd0;
end

always_ff @(posedge clk) begin
	r_idx[0] <= idx_0[13:4];
	r_data[0] <= 64'd0 | (data_0 << ({idx_0[3:0], 2'd0}));
	r_idx[1] <= idx_1[13:4];
	r_data[1] <= 64'd0 | (data_1 << ({idx_1[3:0], 2'd0}));
	r_idx[2] <= idx_2[13:4];
	r_data[2] <= 64'd0 | (data_2 << ({idx_2[3:0], 2'd0}));
	r_idx[3] <= idx_3[13:4];
	r_data[3] <= 64'd0 | (data_3 << ({idx_3[3:0], 2'd0}));
	r_idx[4] <= idx_4[13:4];
	r_data[4] <= 64'd0 | (data_4 << ({idx_4[3:0], 2'd0}));
	r_idx[5] <= idx_5[13:4];
	r_data[5] <= 64'd0 | (data_5 << ({idx_5[3:0], 2'd0}));
	r_idx[6] <= idx_6[13:4];
	r_data[6] <= 64'd0 | (data_6 << ({idx_6[3:0], 2'd0}));
	r_idx[7] <= idx_7[13:4];
	r_data[7] <= 64'd0 | (data_7 << ({idx_7[3:0], 2'd0}));
end

always_comb begin
	busy_out = busy;
end

always_ff @(posedge clk) begin

	if (r_last[2]) begin
		busy <= 1'd1;
		out_cnt <= 10'd0;
	end
	else if (out_cnt == 10'd1023) begin
		busy <= 1'd0;
		out_cnt <= 10'd0;
	end
	else if (busy && out_ready) begin
		busy <= 1'd1;
		out_cnt <= out_cnt + 10'd1;
	end
	else begin
		busy <= busy;
		out_cnt <= out_cnt;
	end
	reading_memory <= busy;
	r_last[0] <= last;
	r_valid[0] <= valid;
	r_last[1] <= r_last[0];
	r_last[2] <= r_last[1];
	r_valid[1] <= r_valid[0];
	r_valid[2] <= r_valid[1];
	r2_idx[0] <= r_idx[0];
	r2_idx[1] <= r_idx[1];
	r2_idx[2] <= r_idx[2];
	r2_idx[3] <= r_idx[3];
	r2_idx[4] <= r_idx[4];
	r2_idx[5] <= r_idx[5];
	r2_idx[6] <= r_idx[6];
	r2_idx[7] <= r_idx[7];
	r3_idx[0] <= r2_idx[0];
	r3_idx[1] <= r2_idx[1];
	r3_idx[2] <= r2_idx[2];
	r3_idx[3] <= r2_idx[3];
	r3_idx[4] <= r2_idx[4];
	r3_idx[5] <= r2_idx[5];
	r3_idx[6] <= r2_idx[6];
	r3_idx[7] <= r2_idx[7];
	r2_data[0] <= r_data[0];
	r2_data[1] <= r_data[1];
	r2_data[2] <= r_data[2];
	r2_data[3] <= r_data[3];
	r2_data[4] <= r_data[4];
	r2_data[5] <= r_data[5];
	r2_data[6] <= r_data[6];
	r2_data[7] <= r_data[7];
	r3_data[0] <= r2_data[0];
	r3_data[1] <= r2_data[1];
	r3_data[2] <= r2_data[2];
	r3_data[3] <= r2_data[3];
	r3_data[4] <= r2_data[4];
	r3_data[5] <= r2_data[5];
	r3_data[6] <= r2_data[6];
	r3_data[7] <= r2_data[7];

	if (busy) begin
		mem_rd_addr[0] <= out_cnt;
		mem_wr_addr[0] <= out_cnt;
		mem_rd_addr[1] <= out_cnt;
		mem_wr_addr[1] <= out_cnt;
		mem_rd_addr[2] <= out_cnt;
		mem_wr_addr[2] <= out_cnt;
		mem_rd_addr[3] <= out_cnt;
		mem_wr_addr[3] <= out_cnt;
		mem_rd_addr[4] <= out_cnt;
		mem_wr_addr[4] <= out_cnt;
		mem_rd_addr[5] <= out_cnt;
		mem_wr_addr[5] <= out_cnt;
		mem_rd_addr[6] <= out_cnt;
		mem_wr_addr[6] <= out_cnt;
		mem_rd_addr[7] <= out_cnt;
		mem_wr_addr[7] <= out_cnt;
	end
	else begin
		mem_rd_addr[0] <= idx_0[13:4];
		mem_wr_addr[0] <= r2_idx[0];
		mem_rd_addr[1] <= idx_1[13:4];
		mem_wr_addr[1] <= r2_idx[1];
		mem_rd_addr[2] <= idx_2[13:4];
		mem_wr_addr[2] <= r2_idx[2];
		mem_rd_addr[3] <= idx_3[13:4];
		mem_wr_addr[3] <= r2_idx[3];
		mem_rd_addr[4] <= idx_4[13:4];
		mem_wr_addr[4] <= r2_idx[4];
		mem_rd_addr[5] <= idx_5[13:4];
		mem_wr_addr[5] <= r2_idx[5];
		mem_rd_addr[6] <= idx_6[13:4];
		mem_wr_addr[6] <= r2_idx[6];
		mem_rd_addr[7] <= idx_7[13:4];
		mem_wr_addr[7] <= r2_idx[7];
	end

	if (r_valid[2][0] || reading_memory) begin
		mem_0[mem_wr_addr[0]] <= in_mem[0];
	end

	if (r_valid[2][1] || reading_memory) begin
		mem_1[mem_wr_addr[1]] <= in_mem[1];
	end

	if (r_valid[2][2] || reading_memory) begin
		mem_2[mem_wr_addr[2]] <= in_mem[2];
	end

	if (r_valid[2][3] || reading_memory) begin
		mem_3[mem_wr_addr[3]] <= in_mem[3];
	end

	if (r_valid[2][4] || reading_memory) begin
		mem_4[mem_wr_addr[4]] <= in_mem[4];
	end

	if (r_valid[2][5] || reading_memory) begin
		mem_5[mem_wr_addr[5]] <= in_mem[5];
	end

	if (r_valid[2][6] || reading_memory) begin
		mem_6[mem_wr_addr[6]] <= in_mem[6];
	end

	if (r_valid[2][7] || reading_memory) begin
		mem_7[mem_wr_addr[7]] <= in_mem[7];
	end
	out_mem[0] <= mem_0[mem_rd_addr[0]];
	out_mem[1] <= mem_1[mem_rd_addr[1]];
	out_mem[2] <= mem_2[mem_rd_addr[2]];
	out_mem[3] <= mem_3[mem_rd_addr[3]];
	out_mem[4] <= mem_4[mem_rd_addr[4]];
	out_mem[5] <= mem_5[mem_rd_addr[5]];
	out_mem[6] <= mem_6[mem_rd_addr[6]];
	out_mem[7] <= mem_7[mem_rd_addr[7]];

	if (busy) begin
		in_mem[0] <= 64'd0;
	end
	else if (r2_idx[0] == r3_idx[0]) begin

		if (r2_data[0][3:0] > in_mem[0][3:0]) begin
			in_mem[0][3:0] <= r2_data[0][3:0];
		end
		else begin
			in_mem[0][3:0] <= in_mem[0][3:0];
		end

		if (r2_data[0][7:4] > in_mem[0][7:4]) begin
			in_mem[0][7:4] <= r2_data[0][7:4];
		end
		else begin
			in_mem[0][7:4] <= in_mem[0][7:4];
		end

		if (r2_data[0][11:8] > in_mem[0][11:8]) begin
			in_mem[0][11:8] <= r2_data[0][11:8];
		end
		else begin
			in_mem[0][11:8] <= in_mem[0][11:8];
		end

		if (r2_data[0][15:12] > in_mem[0][15:12]) begin
			in_mem[0][15:12] <= r2_data[0][15:12];
		end
		else begin
			in_mem[0][15:12] <= in_mem[0][15:12];
		end

		if (r2_data[0][19:16] > in_mem[0][19:16]) begin
			in_mem[0][19:16] <= r2_data[0][19:16];
		end
		else begin
			in_mem[0][19:16] <= in_mem[0][19:16];
		end

		if (r2_data[0][23:20] > in_mem[0][23:20]) begin
			in_mem[0][23:20] <= r2_data[0][23:20];
		end
		else begin
			in_mem[0][23:20] <= in_mem[0][23:20];
		end

		if (r2_data[0][27:24] > in_mem[0][27:24]) begin
			in_mem[0][27:24] <= r2_data[0][27:24];
		end
		else begin
			in_mem[0][27:24] <= in_mem[0][27:24];
		end

		if (r2_data[0][31:28] > in_mem[0][31:28]) begin
			in_mem[0][31:28] <= r2_data[0][31:28];
		end
		else begin
			in_mem[0][31:28] <= in_mem[0][31:28];
		end

		if (r2_data[0][35:32] > in_mem[0][35:32]) begin
			in_mem[0][35:32] <= r2_data[0][35:32];
		end
		else begin
			in_mem[0][35:32] <= in_mem[0][35:32];
		end

		if (r2_data[0][39:36] > in_mem[0][39:36]) begin
			in_mem[0][39:36] <= r2_data[0][39:36];
		end
		else begin
			in_mem[0][39:36] <= in_mem[0][39:36];
		end

		if (r2_data[0][43:40] > in_mem[0][43:40]) begin
			in_mem[0][43:40] <= r2_data[0][43:40];
		end
		else begin
			in_mem[0][43:40] <= in_mem[0][43:40];
		end

		if (r2_data[0][47:44] > in_mem[0][47:44]) begin
			in_mem[0][47:44] <= r2_data[0][47:44];
		end
		else begin
			in_mem[0][47:44] <= in_mem[0][47:44];
		end

		if (r2_data[0][51:48] > in_mem[0][51:48]) begin
			in_mem[0][51:48] <= r2_data[0][51:48];
		end
		else begin
			in_mem[0][51:48] <= in_mem[0][51:48];
		end

		if (r2_data[0][55:52] > in_mem[0][55:52]) begin
			in_mem[0][55:52] <= r2_data[0][55:52];
		end
		else begin
			in_mem[0][55:52] <= in_mem[0][55:52];
		end

		if (r2_data[0][59:56] > in_mem[0][59:56]) begin
			in_mem[0][59:56] <= r2_data[0][59:56];
		end
		else begin
			in_mem[0][59:56] <= in_mem[0][59:56];
		end

		if (r2_data[0][63:60] > in_mem[0][63:60]) begin
			in_mem[0][63:60] <= r2_data[0][63:60];
		end
		else begin
			in_mem[0][63:60] <= in_mem[0][63:60];
		end
	end
	else begin

		if (r2_data[0][3:0] > out_mem[0][3:0]) begin
			in_mem[0][3:0] <= r2_data[0][3:0];
		end
		else begin
			in_mem[0][3:0] <= out_mem[0][3:0];
		end

		if (r2_data[0][7:4] > out_mem[0][7:4]) begin
			in_mem[0][7:4] <= r2_data[0][7:4];
		end
		else begin
			in_mem[0][7:4] <= out_mem[0][7:4];
		end

		if (r2_data[0][11:8] > out_mem[0][11:8]) begin
			in_mem[0][11:8] <= r2_data[0][11:8];
		end
		else begin
			in_mem[0][11:8] <= out_mem[0][11:8];
		end

		if (r2_data[0][15:12] > out_mem[0][15:12]) begin
			in_mem[0][15:12] <= r2_data[0][15:12];
		end
		else begin
			in_mem[0][15:12] <= out_mem[0][15:12];
		end

		if (r2_data[0][19:16] > out_mem[0][19:16]) begin
			in_mem[0][19:16] <= r2_data[0][19:16];
		end
		else begin
			in_mem[0][19:16] <= out_mem[0][19:16];
		end

		if (r2_data[0][23:20] > out_mem[0][23:20]) begin
			in_mem[0][23:20] <= r2_data[0][23:20];
		end
		else begin
			in_mem[0][23:20] <= out_mem[0][23:20];
		end

		if (r2_data[0][27:24] > out_mem[0][27:24]) begin
			in_mem[0][27:24] <= r2_data[0][27:24];
		end
		else begin
			in_mem[0][27:24] <= out_mem[0][27:24];
		end

		if (r2_data[0][31:28] > out_mem[0][31:28]) begin
			in_mem[0][31:28] <= r2_data[0][31:28];
		end
		else begin
			in_mem[0][31:28] <= out_mem[0][31:28];
		end

		if (r2_data[0][35:32] > out_mem[0][35:32]) begin
			in_mem[0][35:32] <= r2_data[0][35:32];
		end
		else begin
			in_mem[0][35:32] <= out_mem[0][35:32];
		end

		if (r2_data[0][39:36] > out_mem[0][39:36]) begin
			in_mem[0][39:36] <= r2_data[0][39:36];
		end
		else begin
			in_mem[0][39:36] <= out_mem[0][39:36];
		end

		if (r2_data[0][43:40] > out_mem[0][43:40]) begin
			in_mem[0][43:40] <= r2_data[0][43:40];
		end
		else begin
			in_mem[0][43:40] <= out_mem[0][43:40];
		end

		if (r2_data[0][47:44] > out_mem[0][47:44]) begin
			in_mem[0][47:44] <= r2_data[0][47:44];
		end
		else begin
			in_mem[0][47:44] <= out_mem[0][47:44];
		end

		if (r2_data[0][51:48] > out_mem[0][51:48]) begin
			in_mem[0][51:48] <= r2_data[0][51:48];
		end
		else begin
			in_mem[0][51:48] <= out_mem[0][51:48];
		end

		if (r2_data[0][55:52] > out_mem[0][55:52]) begin
			in_mem[0][55:52] <= r2_data[0][55:52];
		end
		else begin
			in_mem[0][55:52] <= out_mem[0][55:52];
		end

		if (r2_data[0][59:56] > out_mem[0][59:56]) begin
			in_mem[0][59:56] <= r2_data[0][59:56];
		end
		else begin
			in_mem[0][59:56] <= out_mem[0][59:56];
		end

		if (r2_data[0][63:60] > out_mem[0][63:60]) begin
			in_mem[0][63:60] <= r2_data[0][63:60];
		end
		else begin
			in_mem[0][63:60] <= out_mem[0][63:60];
		end
	end

	if (busy) begin
		in_mem[1] <= 64'd0;
	end
	else if (r2_idx[1] == r3_idx[1]) begin

		if (r2_data[1][3:0] > in_mem[1][3:0]) begin
			in_mem[1][3:0] <= r2_data[1][3:0];
		end
		else begin
			in_mem[1][3:0] <= in_mem[1][3:0];
		end

		if (r2_data[1][7:4] > in_mem[1][7:4]) begin
			in_mem[1][7:4] <= r2_data[1][7:4];
		end
		else begin
			in_mem[1][7:4] <= in_mem[1][7:4];
		end

		if (r2_data[1][11:8] > in_mem[1][11:8]) begin
			in_mem[1][11:8] <= r2_data[1][11:8];
		end
		else begin
			in_mem[1][11:8] <= in_mem[1][11:8];
		end

		if (r2_data[1][15:12] > in_mem[1][15:12]) begin
			in_mem[1][15:12] <= r2_data[1][15:12];
		end
		else begin
			in_mem[1][15:12] <= in_mem[1][15:12];
		end

		if (r2_data[1][19:16] > in_mem[1][19:16]) begin
			in_mem[1][19:16] <= r2_data[1][19:16];
		end
		else begin
			in_mem[1][19:16] <= in_mem[1][19:16];
		end

		if (r2_data[1][23:20] > in_mem[1][23:20]) begin
			in_mem[1][23:20] <= r2_data[1][23:20];
		end
		else begin
			in_mem[1][23:20] <= in_mem[1][23:20];
		end

		if (r2_data[1][27:24] > in_mem[1][27:24]) begin
			in_mem[1][27:24] <= r2_data[1][27:24];
		end
		else begin
			in_mem[1][27:24] <= in_mem[1][27:24];
		end

		if (r2_data[1][31:28] > in_mem[1][31:28]) begin
			in_mem[1][31:28] <= r2_data[1][31:28];
		end
		else begin
			in_mem[1][31:28] <= in_mem[1][31:28];
		end

		if (r2_data[1][35:32] > in_mem[1][35:32]) begin
			in_mem[1][35:32] <= r2_data[1][35:32];
		end
		else begin
			in_mem[1][35:32] <= in_mem[1][35:32];
		end

		if (r2_data[1][39:36] > in_mem[1][39:36]) begin
			in_mem[1][39:36] <= r2_data[1][39:36];
		end
		else begin
			in_mem[1][39:36] <= in_mem[1][39:36];
		end

		if (r2_data[1][43:40] > in_mem[1][43:40]) begin
			in_mem[1][43:40] <= r2_data[1][43:40];
		end
		else begin
			in_mem[1][43:40] <= in_mem[1][43:40];
		end

		if (r2_data[1][47:44] > in_mem[1][47:44]) begin
			in_mem[1][47:44] <= r2_data[1][47:44];
		end
		else begin
			in_mem[1][47:44] <= in_mem[1][47:44];
		end

		if (r2_data[1][51:48] > in_mem[1][51:48]) begin
			in_mem[1][51:48] <= r2_data[1][51:48];
		end
		else begin
			in_mem[1][51:48] <= in_mem[1][51:48];
		end

		if (r2_data[1][55:52] > in_mem[1][55:52]) begin
			in_mem[1][55:52] <= r2_data[1][55:52];
		end
		else begin
			in_mem[1][55:52] <= in_mem[1][55:52];
		end

		if (r2_data[1][59:56] > in_mem[1][59:56]) begin
			in_mem[1][59:56] <= r2_data[1][59:56];
		end
		else begin
			in_mem[1][59:56] <= in_mem[1][59:56];
		end

		if (r2_data[1][63:60] > in_mem[1][63:60]) begin
			in_mem[1][63:60] <= r2_data[1][63:60];
		end
		else begin
			in_mem[1][63:60] <= in_mem[1][63:60];
		end
	end
	else begin

		if (r2_data[1][3:0] > out_mem[1][3:0]) begin
			in_mem[1][3:0] <= r2_data[1][3:0];
		end
		else begin
			in_mem[1][3:0] <= out_mem[1][3:0];
		end

		if (r2_data[1][7:4] > out_mem[1][7:4]) begin
			in_mem[1][7:4] <= r2_data[1][7:4];
		end
		else begin
			in_mem[1][7:4] <= out_mem[1][7:4];
		end

		if (r2_data[1][11:8] > out_mem[1][11:8]) begin
			in_mem[1][11:8] <= r2_data[1][11:8];
		end
		else begin
			in_mem[1][11:8] <= out_mem[1][11:8];
		end

		if (r2_data[1][15:12] > out_mem[1][15:12]) begin
			in_mem[1][15:12] <= r2_data[1][15:12];
		end
		else begin
			in_mem[1][15:12] <= out_mem[1][15:12];
		end

		if (r2_data[1][19:16] > out_mem[1][19:16]) begin
			in_mem[1][19:16] <= r2_data[1][19:16];
		end
		else begin
			in_mem[1][19:16] <= out_mem[1][19:16];
		end

		if (r2_data[1][23:20] > out_mem[1][23:20]) begin
			in_mem[1][23:20] <= r2_data[1][23:20];
		end
		else begin
			in_mem[1][23:20] <= out_mem[1][23:20];
		end

		if (r2_data[1][27:24] > out_mem[1][27:24]) begin
			in_mem[1][27:24] <= r2_data[1][27:24];
		end
		else begin
			in_mem[1][27:24] <= out_mem[1][27:24];
		end

		if (r2_data[1][31:28] > out_mem[1][31:28]) begin
			in_mem[1][31:28] <= r2_data[1][31:28];
		end
		else begin
			in_mem[1][31:28] <= out_mem[1][31:28];
		end

		if (r2_data[1][35:32] > out_mem[1][35:32]) begin
			in_mem[1][35:32] <= r2_data[1][35:32];
		end
		else begin
			in_mem[1][35:32] <= out_mem[1][35:32];
		end

		if (r2_data[1][39:36] > out_mem[1][39:36]) begin
			in_mem[1][39:36] <= r2_data[1][39:36];
		end
		else begin
			in_mem[1][39:36] <= out_mem[1][39:36];
		end

		if (r2_data[1][43:40] > out_mem[1][43:40]) begin
			in_mem[1][43:40] <= r2_data[1][43:40];
		end
		else begin
			in_mem[1][43:40] <= out_mem[1][43:40];
		end

		if (r2_data[1][47:44] > out_mem[1][47:44]) begin
			in_mem[1][47:44] <= r2_data[1][47:44];
		end
		else begin
			in_mem[1][47:44] <= out_mem[1][47:44];
		end

		if (r2_data[1][51:48] > out_mem[1][51:48]) begin
			in_mem[1][51:48] <= r2_data[1][51:48];
		end
		else begin
			in_mem[1][51:48] <= out_mem[1][51:48];
		end

		if (r2_data[1][55:52] > out_mem[1][55:52]) begin
			in_mem[1][55:52] <= r2_data[1][55:52];
		end
		else begin
			in_mem[1][55:52] <= out_mem[1][55:52];
		end

		if (r2_data[1][59:56] > out_mem[1][59:56]) begin
			in_mem[1][59:56] <= r2_data[1][59:56];
		end
		else begin
			in_mem[1][59:56] <= out_mem[1][59:56];
		end

		if (r2_data[1][63:60] > out_mem[1][63:60]) begin
			in_mem[1][63:60] <= r2_data[1][63:60];
		end
		else begin
			in_mem[1][63:60] <= out_mem[1][63:60];
		end
	end

	if (busy) begin
		in_mem[2] <= 64'd0;
	end
	else if (r2_idx[2] == r3_idx[2]) begin

		if (r2_data[2][3:0] > in_mem[2][3:0]) begin
			in_mem[2][3:0] <= r2_data[2][3:0];
		end
		else begin
			in_mem[2][3:0] <= in_mem[2][3:0];
		end

		if (r2_data[2][7:4] > in_mem[2][7:4]) begin
			in_mem[2][7:4] <= r2_data[2][7:4];
		end
		else begin
			in_mem[2][7:4] <= in_mem[2][7:4];
		end

		if (r2_data[2][11:8] > in_mem[2][11:8]) begin
			in_mem[2][11:8] <= r2_data[2][11:8];
		end
		else begin
			in_mem[2][11:8] <= in_mem[2][11:8];
		end

		if (r2_data[2][15:12] > in_mem[2][15:12]) begin
			in_mem[2][15:12] <= r2_data[2][15:12];
		end
		else begin
			in_mem[2][15:12] <= in_mem[2][15:12];
		end

		if (r2_data[2][19:16] > in_mem[2][19:16]) begin
			in_mem[2][19:16] <= r2_data[2][19:16];
		end
		else begin
			in_mem[2][19:16] <= in_mem[2][19:16];
		end

		if (r2_data[2][23:20] > in_mem[2][23:20]) begin
			in_mem[2][23:20] <= r2_data[2][23:20];
		end
		else begin
			in_mem[2][23:20] <= in_mem[2][23:20];
		end

		if (r2_data[2][27:24] > in_mem[2][27:24]) begin
			in_mem[2][27:24] <= r2_data[2][27:24];
		end
		else begin
			in_mem[2][27:24] <= in_mem[2][27:24];
		end

		if (r2_data[2][31:28] > in_mem[2][31:28]) begin
			in_mem[2][31:28] <= r2_data[2][31:28];
		end
		else begin
			in_mem[2][31:28] <= in_mem[2][31:28];
		end

		if (r2_data[2][35:32] > in_mem[2][35:32]) begin
			in_mem[2][35:32] <= r2_data[2][35:32];
		end
		else begin
			in_mem[2][35:32] <= in_mem[2][35:32];
		end

		if (r2_data[2][39:36] > in_mem[2][39:36]) begin
			in_mem[2][39:36] <= r2_data[2][39:36];
		end
		else begin
			in_mem[2][39:36] <= in_mem[2][39:36];
		end

		if (r2_data[2][43:40] > in_mem[2][43:40]) begin
			in_mem[2][43:40] <= r2_data[2][43:40];
		end
		else begin
			in_mem[2][43:40] <= in_mem[2][43:40];
		end

		if (r2_data[2][47:44] > in_mem[2][47:44]) begin
			in_mem[2][47:44] <= r2_data[2][47:44];
		end
		else begin
			in_mem[2][47:44] <= in_mem[2][47:44];
		end

		if (r2_data[2][51:48] > in_mem[2][51:48]) begin
			in_mem[2][51:48] <= r2_data[2][51:48];
		end
		else begin
			in_mem[2][51:48] <= in_mem[2][51:48];
		end

		if (r2_data[2][55:52] > in_mem[2][55:52]) begin
			in_mem[2][55:52] <= r2_data[2][55:52];
		end
		else begin
			in_mem[2][55:52] <= in_mem[2][55:52];
		end

		if (r2_data[2][59:56] > in_mem[2][59:56]) begin
			in_mem[2][59:56] <= r2_data[2][59:56];
		end
		else begin
			in_mem[2][59:56] <= in_mem[2][59:56];
		end

		if (r2_data[2][63:60] > in_mem[2][63:60]) begin
			in_mem[2][63:60] <= r2_data[2][63:60];
		end
		else begin
			in_mem[2][63:60] <= in_mem[2][63:60];
		end
	end
	else begin

		if (r2_data[2][3:0] > out_mem[2][3:0]) begin
			in_mem[2][3:0] <= r2_data[2][3:0];
		end
		else begin
			in_mem[2][3:0] <= out_mem[2][3:0];
		end

		if (r2_data[2][7:4] > out_mem[2][7:4]) begin
			in_mem[2][7:4] <= r2_data[2][7:4];
		end
		else begin
			in_mem[2][7:4] <= out_mem[2][7:4];
		end

		if (r2_data[2][11:8] > out_mem[2][11:8]) begin
			in_mem[2][11:8] <= r2_data[2][11:8];
		end
		else begin
			in_mem[2][11:8] <= out_mem[2][11:8];
		end

		if (r2_data[2][15:12] > out_mem[2][15:12]) begin
			in_mem[2][15:12] <= r2_data[2][15:12];
		end
		else begin
			in_mem[2][15:12] <= out_mem[2][15:12];
		end

		if (r2_data[2][19:16] > out_mem[2][19:16]) begin
			in_mem[2][19:16] <= r2_data[2][19:16];
		end
		else begin
			in_mem[2][19:16] <= out_mem[2][19:16];
		end

		if (r2_data[2][23:20] > out_mem[2][23:20]) begin
			in_mem[2][23:20] <= r2_data[2][23:20];
		end
		else begin
			in_mem[2][23:20] <= out_mem[2][23:20];
		end

		if (r2_data[2][27:24] > out_mem[2][27:24]) begin
			in_mem[2][27:24] <= r2_data[2][27:24];
		end
		else begin
			in_mem[2][27:24] <= out_mem[2][27:24];
		end

		if (r2_data[2][31:28] > out_mem[2][31:28]) begin
			in_mem[2][31:28] <= r2_data[2][31:28];
		end
		else begin
			in_mem[2][31:28] <= out_mem[2][31:28];
		end

		if (r2_data[2][35:32] > out_mem[2][35:32]) begin
			in_mem[2][35:32] <= r2_data[2][35:32];
		end
		else begin
			in_mem[2][35:32] <= out_mem[2][35:32];
		end

		if (r2_data[2][39:36] > out_mem[2][39:36]) begin
			in_mem[2][39:36] <= r2_data[2][39:36];
		end
		else begin
			in_mem[2][39:36] <= out_mem[2][39:36];
		end

		if (r2_data[2][43:40] > out_mem[2][43:40]) begin
			in_mem[2][43:40] <= r2_data[2][43:40];
		end
		else begin
			in_mem[2][43:40] <= out_mem[2][43:40];
		end

		if (r2_data[2][47:44] > out_mem[2][47:44]) begin
			in_mem[2][47:44] <= r2_data[2][47:44];
		end
		else begin
			in_mem[2][47:44] <= out_mem[2][47:44];
		end

		if (r2_data[2][51:48] > out_mem[2][51:48]) begin
			in_mem[2][51:48] <= r2_data[2][51:48];
		end
		else begin
			in_mem[2][51:48] <= out_mem[2][51:48];
		end

		if (r2_data[2][55:52] > out_mem[2][55:52]) begin
			in_mem[2][55:52] <= r2_data[2][55:52];
		end
		else begin
			in_mem[2][55:52] <= out_mem[2][55:52];
		end

		if (r2_data[2][59:56] > out_mem[2][59:56]) begin
			in_mem[2][59:56] <= r2_data[2][59:56];
		end
		else begin
			in_mem[2][59:56] <= out_mem[2][59:56];
		end

		if (r2_data[2][63:60] > out_mem[2][63:60]) begin
			in_mem[2][63:60] <= r2_data[2][63:60];
		end
		else begin
			in_mem[2][63:60] <= out_mem[2][63:60];
		end
	end

	if (busy) begin
		in_mem[3] <= 64'd0;
	end
	else if (r2_idx[3] == r3_idx[3]) begin

		if (r2_data[3][3:0] > in_mem[3][3:0]) begin
			in_mem[3][3:0] <= r2_data[3][3:0];
		end
		else begin
			in_mem[3][3:0] <= in_mem[3][3:0];
		end

		if (r2_data[3][7:4] > in_mem[3][7:4]) begin
			in_mem[3][7:4] <= r2_data[3][7:4];
		end
		else begin
			in_mem[3][7:4] <= in_mem[3][7:4];
		end

		if (r2_data[3][11:8] > in_mem[3][11:8]) begin
			in_mem[3][11:8] <= r2_data[3][11:8];
		end
		else begin
			in_mem[3][11:8] <= in_mem[3][11:8];
		end

		if (r2_data[3][15:12] > in_mem[3][15:12]) begin
			in_mem[3][15:12] <= r2_data[3][15:12];
		end
		else begin
			in_mem[3][15:12] <= in_mem[3][15:12];
		end

		if (r2_data[3][19:16] > in_mem[3][19:16]) begin
			in_mem[3][19:16] <= r2_data[3][19:16];
		end
		else begin
			in_mem[3][19:16] <= in_mem[3][19:16];
		end

		if (r2_data[3][23:20] > in_mem[3][23:20]) begin
			in_mem[3][23:20] <= r2_data[3][23:20];
		end
		else begin
			in_mem[3][23:20] <= in_mem[3][23:20];
		end

		if (r2_data[3][27:24] > in_mem[3][27:24]) begin
			in_mem[3][27:24] <= r2_data[3][27:24];
		end
		else begin
			in_mem[3][27:24] <= in_mem[3][27:24];
		end

		if (r2_data[3][31:28] > in_mem[3][31:28]) begin
			in_mem[3][31:28] <= r2_data[3][31:28];
		end
		else begin
			in_mem[3][31:28] <= in_mem[3][31:28];
		end

		if (r2_data[3][35:32] > in_mem[3][35:32]) begin
			in_mem[3][35:32] <= r2_data[3][35:32];
		end
		else begin
			in_mem[3][35:32] <= in_mem[3][35:32];
		end

		if (r2_data[3][39:36] > in_mem[3][39:36]) begin
			in_mem[3][39:36] <= r2_data[3][39:36];
		end
		else begin
			in_mem[3][39:36] <= in_mem[3][39:36];
		end

		if (r2_data[3][43:40] > in_mem[3][43:40]) begin
			in_mem[3][43:40] <= r2_data[3][43:40];
		end
		else begin
			in_mem[3][43:40] <= in_mem[3][43:40];
		end

		if (r2_data[3][47:44] > in_mem[3][47:44]) begin
			in_mem[3][47:44] <= r2_data[3][47:44];
		end
		else begin
			in_mem[3][47:44] <= in_mem[3][47:44];
		end

		if (r2_data[3][51:48] > in_mem[3][51:48]) begin
			in_mem[3][51:48] <= r2_data[3][51:48];
		end
		else begin
			in_mem[3][51:48] <= in_mem[3][51:48];
		end

		if (r2_data[3][55:52] > in_mem[3][55:52]) begin
			in_mem[3][55:52] <= r2_data[3][55:52];
		end
		else begin
			in_mem[3][55:52] <= in_mem[3][55:52];
		end

		if (r2_data[3][59:56] > in_mem[3][59:56]) begin
			in_mem[3][59:56] <= r2_data[3][59:56];
		end
		else begin
			in_mem[3][59:56] <= in_mem[3][59:56];
		end

		if (r2_data[3][63:60] > in_mem[3][63:60]) begin
			in_mem[3][63:60] <= r2_data[3][63:60];
		end
		else begin
			in_mem[3][63:60] <= in_mem[3][63:60];
		end
	end
	else begin

		if (r2_data[3][3:0] > out_mem[3][3:0]) begin
			in_mem[3][3:0] <= r2_data[3][3:0];
		end
		else begin
			in_mem[3][3:0] <= out_mem[3][3:0];
		end

		if (r2_data[3][7:4] > out_mem[3][7:4]) begin
			in_mem[3][7:4] <= r2_data[3][7:4];
		end
		else begin
			in_mem[3][7:4] <= out_mem[3][7:4];
		end

		if (r2_data[3][11:8] > out_mem[3][11:8]) begin
			in_mem[3][11:8] <= r2_data[3][11:8];
		end
		else begin
			in_mem[3][11:8] <= out_mem[3][11:8];
		end

		if (r2_data[3][15:12] > out_mem[3][15:12]) begin
			in_mem[3][15:12] <= r2_data[3][15:12];
		end
		else begin
			in_mem[3][15:12] <= out_mem[3][15:12];
		end

		if (r2_data[3][19:16] > out_mem[3][19:16]) begin
			in_mem[3][19:16] <= r2_data[3][19:16];
		end
		else begin
			in_mem[3][19:16] <= out_mem[3][19:16];
		end

		if (r2_data[3][23:20] > out_mem[3][23:20]) begin
			in_mem[3][23:20] <= r2_data[3][23:20];
		end
		else begin
			in_mem[3][23:20] <= out_mem[3][23:20];
		end

		if (r2_data[3][27:24] > out_mem[3][27:24]) begin
			in_mem[3][27:24] <= r2_data[3][27:24];
		end
		else begin
			in_mem[3][27:24] <= out_mem[3][27:24];
		end

		if (r2_data[3][31:28] > out_mem[3][31:28]) begin
			in_mem[3][31:28] <= r2_data[3][31:28];
		end
		else begin
			in_mem[3][31:28] <= out_mem[3][31:28];
		end

		if (r2_data[3][35:32] > out_mem[3][35:32]) begin
			in_mem[3][35:32] <= r2_data[3][35:32];
		end
		else begin
			in_mem[3][35:32] <= out_mem[3][35:32];
		end

		if (r2_data[3][39:36] > out_mem[3][39:36]) begin
			in_mem[3][39:36] <= r2_data[3][39:36];
		end
		else begin
			in_mem[3][39:36] <= out_mem[3][39:36];
		end

		if (r2_data[3][43:40] > out_mem[3][43:40]) begin
			in_mem[3][43:40] <= r2_data[3][43:40];
		end
		else begin
			in_mem[3][43:40] <= out_mem[3][43:40];
		end

		if (r2_data[3][47:44] > out_mem[3][47:44]) begin
			in_mem[3][47:44] <= r2_data[3][47:44];
		end
		else begin
			in_mem[3][47:44] <= out_mem[3][47:44];
		end

		if (r2_data[3][51:48] > out_mem[3][51:48]) begin
			in_mem[3][51:48] <= r2_data[3][51:48];
		end
		else begin
			in_mem[3][51:48] <= out_mem[3][51:48];
		end

		if (r2_data[3][55:52] > out_mem[3][55:52]) begin
			in_mem[3][55:52] <= r2_data[3][55:52];
		end
		else begin
			in_mem[3][55:52] <= out_mem[3][55:52];
		end

		if (r2_data[3][59:56] > out_mem[3][59:56]) begin
			in_mem[3][59:56] <= r2_data[3][59:56];
		end
		else begin
			in_mem[3][59:56] <= out_mem[3][59:56];
		end

		if (r2_data[3][63:60] > out_mem[3][63:60]) begin
			in_mem[3][63:60] <= r2_data[3][63:60];
		end
		else begin
			in_mem[3][63:60] <= out_mem[3][63:60];
		end
	end

	if (busy) begin
		in_mem[4] <= 64'd0;
	end
	else if (r2_idx[4] == r3_idx[4]) begin

		if (r2_data[4][3:0] > in_mem[4][3:0]) begin
			in_mem[4][3:0] <= r2_data[4][3:0];
		end
		else begin
			in_mem[4][3:0] <= in_mem[4][3:0];
		end

		if (r2_data[4][7:4] > in_mem[4][7:4]) begin
			in_mem[4][7:4] <= r2_data[4][7:4];
		end
		else begin
			in_mem[4][7:4] <= in_mem[4][7:4];
		end

		if (r2_data[4][11:8] > in_mem[4][11:8]) begin
			in_mem[4][11:8] <= r2_data[4][11:8];
		end
		else begin
			in_mem[4][11:8] <= in_mem[4][11:8];
		end

		if (r2_data[4][15:12] > in_mem[4][15:12]) begin
			in_mem[4][15:12] <= r2_data[4][15:12];
		end
		else begin
			in_mem[4][15:12] <= in_mem[4][15:12];
		end

		if (r2_data[4][19:16] > in_mem[4][19:16]) begin
			in_mem[4][19:16] <= r2_data[4][19:16];
		end
		else begin
			in_mem[4][19:16] <= in_mem[4][19:16];
		end

		if (r2_data[4][23:20] > in_mem[4][23:20]) begin
			in_mem[4][23:20] <= r2_data[4][23:20];
		end
		else begin
			in_mem[4][23:20] <= in_mem[4][23:20];
		end

		if (r2_data[4][27:24] > in_mem[4][27:24]) begin
			in_mem[4][27:24] <= r2_data[4][27:24];
		end
		else begin
			in_mem[4][27:24] <= in_mem[4][27:24];
		end

		if (r2_data[4][31:28] > in_mem[4][31:28]) begin
			in_mem[4][31:28] <= r2_data[4][31:28];
		end
		else begin
			in_mem[4][31:28] <= in_mem[4][31:28];
		end

		if (r2_data[4][35:32] > in_mem[4][35:32]) begin
			in_mem[4][35:32] <= r2_data[4][35:32];
		end
		else begin
			in_mem[4][35:32] <= in_mem[4][35:32];
		end

		if (r2_data[4][39:36] > in_mem[4][39:36]) begin
			in_mem[4][39:36] <= r2_data[4][39:36];
		end
		else begin
			in_mem[4][39:36] <= in_mem[4][39:36];
		end

		if (r2_data[4][43:40] > in_mem[4][43:40]) begin
			in_mem[4][43:40] <= r2_data[4][43:40];
		end
		else begin
			in_mem[4][43:40] <= in_mem[4][43:40];
		end

		if (r2_data[4][47:44] > in_mem[4][47:44]) begin
			in_mem[4][47:44] <= r2_data[4][47:44];
		end
		else begin
			in_mem[4][47:44] <= in_mem[4][47:44];
		end

		if (r2_data[4][51:48] > in_mem[4][51:48]) begin
			in_mem[4][51:48] <= r2_data[4][51:48];
		end
		else begin
			in_mem[4][51:48] <= in_mem[4][51:48];
		end

		if (r2_data[4][55:52] > in_mem[4][55:52]) begin
			in_mem[4][55:52] <= r2_data[4][55:52];
		end
		else begin
			in_mem[4][55:52] <= in_mem[4][55:52];
		end

		if (r2_data[4][59:56] > in_mem[4][59:56]) begin
			in_mem[4][59:56] <= r2_data[4][59:56];
		end
		else begin
			in_mem[4][59:56] <= in_mem[4][59:56];
		end

		if (r2_data[4][63:60] > in_mem[4][63:60]) begin
			in_mem[4][63:60] <= r2_data[4][63:60];
		end
		else begin
			in_mem[4][63:60] <= in_mem[4][63:60];
		end
	end
	else begin

		if (r2_data[4][3:0] > out_mem[4][3:0]) begin
			in_mem[4][3:0] <= r2_data[4][3:0];
		end
		else begin
			in_mem[4][3:0] <= out_mem[4][3:0];
		end

		if (r2_data[4][7:4] > out_mem[4][7:4]) begin
			in_mem[4][7:4] <= r2_data[4][7:4];
		end
		else begin
			in_mem[4][7:4] <= out_mem[4][7:4];
		end

		if (r2_data[4][11:8] > out_mem[4][11:8]) begin
			in_mem[4][11:8] <= r2_data[4][11:8];
		end
		else begin
			in_mem[4][11:8] <= out_mem[4][11:8];
		end

		if (r2_data[4][15:12] > out_mem[4][15:12]) begin
			in_mem[4][15:12] <= r2_data[4][15:12];
		end
		else begin
			in_mem[4][15:12] <= out_mem[4][15:12];
		end

		if (r2_data[4][19:16] > out_mem[4][19:16]) begin
			in_mem[4][19:16] <= r2_data[4][19:16];
		end
		else begin
			in_mem[4][19:16] <= out_mem[4][19:16];
		end

		if (r2_data[4][23:20] > out_mem[4][23:20]) begin
			in_mem[4][23:20] <= r2_data[4][23:20];
		end
		else begin
			in_mem[4][23:20] <= out_mem[4][23:20];
		end

		if (r2_data[4][27:24] > out_mem[4][27:24]) begin
			in_mem[4][27:24] <= r2_data[4][27:24];
		end
		else begin
			in_mem[4][27:24] <= out_mem[4][27:24];
		end

		if (r2_data[4][31:28] > out_mem[4][31:28]) begin
			in_mem[4][31:28] <= r2_data[4][31:28];
		end
		else begin
			in_mem[4][31:28] <= out_mem[4][31:28];
		end

		if (r2_data[4][35:32] > out_mem[4][35:32]) begin
			in_mem[4][35:32] <= r2_data[4][35:32];
		end
		else begin
			in_mem[4][35:32] <= out_mem[4][35:32];
		end

		if (r2_data[4][39:36] > out_mem[4][39:36]) begin
			in_mem[4][39:36] <= r2_data[4][39:36];
		end
		else begin
			in_mem[4][39:36] <= out_mem[4][39:36];
		end

		if (r2_data[4][43:40] > out_mem[4][43:40]) begin
			in_mem[4][43:40] <= r2_data[4][43:40];
		end
		else begin
			in_mem[4][43:40] <= out_mem[4][43:40];
		end

		if (r2_data[4][47:44] > out_mem[4][47:44]) begin
			in_mem[4][47:44] <= r2_data[4][47:44];
		end
		else begin
			in_mem[4][47:44] <= out_mem[4][47:44];
		end

		if (r2_data[4][51:48] > out_mem[4][51:48]) begin
			in_mem[4][51:48] <= r2_data[4][51:48];
		end
		else begin
			in_mem[4][51:48] <= out_mem[4][51:48];
		end

		if (r2_data[4][55:52] > out_mem[4][55:52]) begin
			in_mem[4][55:52] <= r2_data[4][55:52];
		end
		else begin
			in_mem[4][55:52] <= out_mem[4][55:52];
		end

		if (r2_data[4][59:56] > out_mem[4][59:56]) begin
			in_mem[4][59:56] <= r2_data[4][59:56];
		end
		else begin
			in_mem[4][59:56] <= out_mem[4][59:56];
		end

		if (r2_data[4][63:60] > out_mem[4][63:60]) begin
			in_mem[4][63:60] <= r2_data[4][63:60];
		end
		else begin
			in_mem[4][63:60] <= out_mem[4][63:60];
		end
	end

	if (busy) begin
		in_mem[5] <= 64'd0;
	end
	else if (r2_idx[5] == r3_idx[5]) begin

		if (r2_data[5][3:0] > in_mem[5][3:0]) begin
			in_mem[5][3:0] <= r2_data[5][3:0];
		end
		else begin
			in_mem[5][3:0] <= in_mem[5][3:0];
		end

		if (r2_data[5][7:4] > in_mem[5][7:4]) begin
			in_mem[5][7:4] <= r2_data[5][7:4];
		end
		else begin
			in_mem[5][7:4] <= in_mem[5][7:4];
		end

		if (r2_data[5][11:8] > in_mem[5][11:8]) begin
			in_mem[5][11:8] <= r2_data[5][11:8];
		end
		else begin
			in_mem[5][11:8] <= in_mem[5][11:8];
		end

		if (r2_data[5][15:12] > in_mem[5][15:12]) begin
			in_mem[5][15:12] <= r2_data[5][15:12];
		end
		else begin
			in_mem[5][15:12] <= in_mem[5][15:12];
		end

		if (r2_data[5][19:16] > in_mem[5][19:16]) begin
			in_mem[5][19:16] <= r2_data[5][19:16];
		end
		else begin
			in_mem[5][19:16] <= in_mem[5][19:16];
		end

		if (r2_data[5][23:20] > in_mem[5][23:20]) begin
			in_mem[5][23:20] <= r2_data[5][23:20];
		end
		else begin
			in_mem[5][23:20] <= in_mem[5][23:20];
		end

		if (r2_data[5][27:24] > in_mem[5][27:24]) begin
			in_mem[5][27:24] <= r2_data[5][27:24];
		end
		else begin
			in_mem[5][27:24] <= in_mem[5][27:24];
		end

		if (r2_data[5][31:28] > in_mem[5][31:28]) begin
			in_mem[5][31:28] <= r2_data[5][31:28];
		end
		else begin
			in_mem[5][31:28] <= in_mem[5][31:28];
		end

		if (r2_data[5][35:32] > in_mem[5][35:32]) begin
			in_mem[5][35:32] <= r2_data[5][35:32];
		end
		else begin
			in_mem[5][35:32] <= in_mem[5][35:32];
		end

		if (r2_data[5][39:36] > in_mem[5][39:36]) begin
			in_mem[5][39:36] <= r2_data[5][39:36];
		end
		else begin
			in_mem[5][39:36] <= in_mem[5][39:36];
		end

		if (r2_data[5][43:40] > in_mem[5][43:40]) begin
			in_mem[5][43:40] <= r2_data[5][43:40];
		end
		else begin
			in_mem[5][43:40] <= in_mem[5][43:40];
		end

		if (r2_data[5][47:44] > in_mem[5][47:44]) begin
			in_mem[5][47:44] <= r2_data[5][47:44];
		end
		else begin
			in_mem[5][47:44] <= in_mem[5][47:44];
		end

		if (r2_data[5][51:48] > in_mem[5][51:48]) begin
			in_mem[5][51:48] <= r2_data[5][51:48];
		end
		else begin
			in_mem[5][51:48] <= in_mem[5][51:48];
		end

		if (r2_data[5][55:52] > in_mem[5][55:52]) begin
			in_mem[5][55:52] <= r2_data[5][55:52];
		end
		else begin
			in_mem[5][55:52] <= in_mem[5][55:52];
		end

		if (r2_data[5][59:56] > in_mem[5][59:56]) begin
			in_mem[5][59:56] <= r2_data[5][59:56];
		end
		else begin
			in_mem[5][59:56] <= in_mem[5][59:56];
		end

		if (r2_data[5][63:60] > in_mem[5][63:60]) begin
			in_mem[5][63:60] <= r2_data[5][63:60];
		end
		else begin
			in_mem[5][63:60] <= in_mem[5][63:60];
		end
	end
	else begin

		if (r2_data[5][3:0] > out_mem[5][3:0]) begin
			in_mem[5][3:0] <= r2_data[5][3:0];
		end
		else begin
			in_mem[5][3:0] <= out_mem[5][3:0];
		end

		if (r2_data[5][7:4] > out_mem[5][7:4]) begin
			in_mem[5][7:4] <= r2_data[5][7:4];
		end
		else begin
			in_mem[5][7:4] <= out_mem[5][7:4];
		end

		if (r2_data[5][11:8] > out_mem[5][11:8]) begin
			in_mem[5][11:8] <= r2_data[5][11:8];
		end
		else begin
			in_mem[5][11:8] <= out_mem[5][11:8];
		end

		if (r2_data[5][15:12] > out_mem[5][15:12]) begin
			in_mem[5][15:12] <= r2_data[5][15:12];
		end
		else begin
			in_mem[5][15:12] <= out_mem[5][15:12];
		end

		if (r2_data[5][19:16] > out_mem[5][19:16]) begin
			in_mem[5][19:16] <= r2_data[5][19:16];
		end
		else begin
			in_mem[5][19:16] <= out_mem[5][19:16];
		end

		if (r2_data[5][23:20] > out_mem[5][23:20]) begin
			in_mem[5][23:20] <= r2_data[5][23:20];
		end
		else begin
			in_mem[5][23:20] <= out_mem[5][23:20];
		end

		if (r2_data[5][27:24] > out_mem[5][27:24]) begin
			in_mem[5][27:24] <= r2_data[5][27:24];
		end
		else begin
			in_mem[5][27:24] <= out_mem[5][27:24];
		end

		if (r2_data[5][31:28] > out_mem[5][31:28]) begin
			in_mem[5][31:28] <= r2_data[5][31:28];
		end
		else begin
			in_mem[5][31:28] <= out_mem[5][31:28];
		end

		if (r2_data[5][35:32] > out_mem[5][35:32]) begin
			in_mem[5][35:32] <= r2_data[5][35:32];
		end
		else begin
			in_mem[5][35:32] <= out_mem[5][35:32];
		end

		if (r2_data[5][39:36] > out_mem[5][39:36]) begin
			in_mem[5][39:36] <= r2_data[5][39:36];
		end
		else begin
			in_mem[5][39:36] <= out_mem[5][39:36];
		end

		if (r2_data[5][43:40] > out_mem[5][43:40]) begin
			in_mem[5][43:40] <= r2_data[5][43:40];
		end
		else begin
			in_mem[5][43:40] <= out_mem[5][43:40];
		end

		if (r2_data[5][47:44] > out_mem[5][47:44]) begin
			in_mem[5][47:44] <= r2_data[5][47:44];
		end
		else begin
			in_mem[5][47:44] <= out_mem[5][47:44];
		end

		if (r2_data[5][51:48] > out_mem[5][51:48]) begin
			in_mem[5][51:48] <= r2_data[5][51:48];
		end
		else begin
			in_mem[5][51:48] <= out_mem[5][51:48];
		end

		if (r2_data[5][55:52] > out_mem[5][55:52]) begin
			in_mem[5][55:52] <= r2_data[5][55:52];
		end
		else begin
			in_mem[5][55:52] <= out_mem[5][55:52];
		end

		if (r2_data[5][59:56] > out_mem[5][59:56]) begin
			in_mem[5][59:56] <= r2_data[5][59:56];
		end
		else begin
			in_mem[5][59:56] <= out_mem[5][59:56];
		end

		if (r2_data[5][63:60] > out_mem[5][63:60]) begin
			in_mem[5][63:60] <= r2_data[5][63:60];
		end
		else begin
			in_mem[5][63:60] <= out_mem[5][63:60];
		end
	end

	if (busy) begin
		in_mem[6] <= 64'd0;
	end
	else if (r2_idx[6] == r3_idx[6]) begin

		if (r2_data[6][3:0] > in_mem[6][3:0]) begin
			in_mem[6][3:0] <= r2_data[6][3:0];
		end
		else begin
			in_mem[6][3:0] <= in_mem[6][3:0];
		end

		if (r2_data[6][7:4] > in_mem[6][7:4]) begin
			in_mem[6][7:4] <= r2_data[6][7:4];
		end
		else begin
			in_mem[6][7:4] <= in_mem[6][7:4];
		end

		if (r2_data[6][11:8] > in_mem[6][11:8]) begin
			in_mem[6][11:8] <= r2_data[6][11:8];
		end
		else begin
			in_mem[6][11:8] <= in_mem[6][11:8];
		end

		if (r2_data[6][15:12] > in_mem[6][15:12]) begin
			in_mem[6][15:12] <= r2_data[6][15:12];
		end
		else begin
			in_mem[6][15:12] <= in_mem[6][15:12];
		end

		if (r2_data[6][19:16] > in_mem[6][19:16]) begin
			in_mem[6][19:16] <= r2_data[6][19:16];
		end
		else begin
			in_mem[6][19:16] <= in_mem[6][19:16];
		end

		if (r2_data[6][23:20] > in_mem[6][23:20]) begin
			in_mem[6][23:20] <= r2_data[6][23:20];
		end
		else begin
			in_mem[6][23:20] <= in_mem[6][23:20];
		end

		if (r2_data[6][27:24] > in_mem[6][27:24]) begin
			in_mem[6][27:24] <= r2_data[6][27:24];
		end
		else begin
			in_mem[6][27:24] <= in_mem[6][27:24];
		end

		if (r2_data[6][31:28] > in_mem[6][31:28]) begin
			in_mem[6][31:28] <= r2_data[6][31:28];
		end
		else begin
			in_mem[6][31:28] <= in_mem[6][31:28];
		end

		if (r2_data[6][35:32] > in_mem[6][35:32]) begin
			in_mem[6][35:32] <= r2_data[6][35:32];
		end
		else begin
			in_mem[6][35:32] <= in_mem[6][35:32];
		end

		if (r2_data[6][39:36] > in_mem[6][39:36]) begin
			in_mem[6][39:36] <= r2_data[6][39:36];
		end
		else begin
			in_mem[6][39:36] <= in_mem[6][39:36];
		end

		if (r2_data[6][43:40] > in_mem[6][43:40]) begin
			in_mem[6][43:40] <= r2_data[6][43:40];
		end
		else begin
			in_mem[6][43:40] <= in_mem[6][43:40];
		end

		if (r2_data[6][47:44] > in_mem[6][47:44]) begin
			in_mem[6][47:44] <= r2_data[6][47:44];
		end
		else begin
			in_mem[6][47:44] <= in_mem[6][47:44];
		end

		if (r2_data[6][51:48] > in_mem[6][51:48]) begin
			in_mem[6][51:48] <= r2_data[6][51:48];
		end
		else begin
			in_mem[6][51:48] <= in_mem[6][51:48];
		end

		if (r2_data[6][55:52] > in_mem[6][55:52]) begin
			in_mem[6][55:52] <= r2_data[6][55:52];
		end
		else begin
			in_mem[6][55:52] <= in_mem[6][55:52];
		end

		if (r2_data[6][59:56] > in_mem[6][59:56]) begin
			in_mem[6][59:56] <= r2_data[6][59:56];
		end
		else begin
			in_mem[6][59:56] <= in_mem[6][59:56];
		end

		if (r2_data[6][63:60] > in_mem[6][63:60]) begin
			in_mem[6][63:60] <= r2_data[6][63:60];
		end
		else begin
			in_mem[6][63:60] <= in_mem[6][63:60];
		end
	end
	else begin

		if (r2_data[6][3:0] > out_mem[6][3:0]) begin
			in_mem[6][3:0] <= r2_data[6][3:0];
		end
		else begin
			in_mem[6][3:0] <= out_mem[6][3:0];
		end

		if (r2_data[6][7:4] > out_mem[6][7:4]) begin
			in_mem[6][7:4] <= r2_data[6][7:4];
		end
		else begin
			in_mem[6][7:4] <= out_mem[6][7:4];
		end

		if (r2_data[6][11:8] > out_mem[6][11:8]) begin
			in_mem[6][11:8] <= r2_data[6][11:8];
		end
		else begin
			in_mem[6][11:8] <= out_mem[6][11:8];
		end

		if (r2_data[6][15:12] > out_mem[6][15:12]) begin
			in_mem[6][15:12] <= r2_data[6][15:12];
		end
		else begin
			in_mem[6][15:12] <= out_mem[6][15:12];
		end

		if (r2_data[6][19:16] > out_mem[6][19:16]) begin
			in_mem[6][19:16] <= r2_data[6][19:16];
		end
		else begin
			in_mem[6][19:16] <= out_mem[6][19:16];
		end

		if (r2_data[6][23:20] > out_mem[6][23:20]) begin
			in_mem[6][23:20] <= r2_data[6][23:20];
		end
		else begin
			in_mem[6][23:20] <= out_mem[6][23:20];
		end

		if (r2_data[6][27:24] > out_mem[6][27:24]) begin
			in_mem[6][27:24] <= r2_data[6][27:24];
		end
		else begin
			in_mem[6][27:24] <= out_mem[6][27:24];
		end

		if (r2_data[6][31:28] > out_mem[6][31:28]) begin
			in_mem[6][31:28] <= r2_data[6][31:28];
		end
		else begin
			in_mem[6][31:28] <= out_mem[6][31:28];
		end

		if (r2_data[6][35:32] > out_mem[6][35:32]) begin
			in_mem[6][35:32] <= r2_data[6][35:32];
		end
		else begin
			in_mem[6][35:32] <= out_mem[6][35:32];
		end

		if (r2_data[6][39:36] > out_mem[6][39:36]) begin
			in_mem[6][39:36] <= r2_data[6][39:36];
		end
		else begin
			in_mem[6][39:36] <= out_mem[6][39:36];
		end

		if (r2_data[6][43:40] > out_mem[6][43:40]) begin
			in_mem[6][43:40] <= r2_data[6][43:40];
		end
		else begin
			in_mem[6][43:40] <= out_mem[6][43:40];
		end

		if (r2_data[6][47:44] > out_mem[6][47:44]) begin
			in_mem[6][47:44] <= r2_data[6][47:44];
		end
		else begin
			in_mem[6][47:44] <= out_mem[6][47:44];
		end

		if (r2_data[6][51:48] > out_mem[6][51:48]) begin
			in_mem[6][51:48] <= r2_data[6][51:48];
		end
		else begin
			in_mem[6][51:48] <= out_mem[6][51:48];
		end

		if (r2_data[6][55:52] > out_mem[6][55:52]) begin
			in_mem[6][55:52] <= r2_data[6][55:52];
		end
		else begin
			in_mem[6][55:52] <= out_mem[6][55:52];
		end

		if (r2_data[6][59:56] > out_mem[6][59:56]) begin
			in_mem[6][59:56] <= r2_data[6][59:56];
		end
		else begin
			in_mem[6][59:56] <= out_mem[6][59:56];
		end

		if (r2_data[6][63:60] > out_mem[6][63:60]) begin
			in_mem[6][63:60] <= r2_data[6][63:60];
		end
		else begin
			in_mem[6][63:60] <= out_mem[6][63:60];
		end
	end

	if (busy) begin
		in_mem[7] <= 64'd0;
	end
	else if (r2_idx[7] == r3_idx[7]) begin

		if (r2_data[7][3:0] > in_mem[7][3:0]) begin
			in_mem[7][3:0] <= r2_data[7][3:0];
		end
		else begin
			in_mem[7][3:0] <= in_mem[7][3:0];
		end

		if (r2_data[7][7:4] > in_mem[7][7:4]) begin
			in_mem[7][7:4] <= r2_data[7][7:4];
		end
		else begin
			in_mem[7][7:4] <= in_mem[7][7:4];
		end

		if (r2_data[7][11:8] > in_mem[7][11:8]) begin
			in_mem[7][11:8] <= r2_data[7][11:8];
		end
		else begin
			in_mem[7][11:8] <= in_mem[7][11:8];
		end

		if (r2_data[7][15:12] > in_mem[7][15:12]) begin
			in_mem[7][15:12] <= r2_data[7][15:12];
		end
		else begin
			in_mem[7][15:12] <= in_mem[7][15:12];
		end

		if (r2_data[7][19:16] > in_mem[7][19:16]) begin
			in_mem[7][19:16] <= r2_data[7][19:16];
		end
		else begin
			in_mem[7][19:16] <= in_mem[7][19:16];
		end

		if (r2_data[7][23:20] > in_mem[7][23:20]) begin
			in_mem[7][23:20] <= r2_data[7][23:20];
		end
		else begin
			in_mem[7][23:20] <= in_mem[7][23:20];
		end

		if (r2_data[7][27:24] > in_mem[7][27:24]) begin
			in_mem[7][27:24] <= r2_data[7][27:24];
		end
		else begin
			in_mem[7][27:24] <= in_mem[7][27:24];
		end

		if (r2_data[7][31:28] > in_mem[7][31:28]) begin
			in_mem[7][31:28] <= r2_data[7][31:28];
		end
		else begin
			in_mem[7][31:28] <= in_mem[7][31:28];
		end

		if (r2_data[7][35:32] > in_mem[7][35:32]) begin
			in_mem[7][35:32] <= r2_data[7][35:32];
		end
		else begin
			in_mem[7][35:32] <= in_mem[7][35:32];
		end

		if (r2_data[7][39:36] > in_mem[7][39:36]) begin
			in_mem[7][39:36] <= r2_data[7][39:36];
		end
		else begin
			in_mem[7][39:36] <= in_mem[7][39:36];
		end

		if (r2_data[7][43:40] > in_mem[7][43:40]) begin
			in_mem[7][43:40] <= r2_data[7][43:40];
		end
		else begin
			in_mem[7][43:40] <= in_mem[7][43:40];
		end

		if (r2_data[7][47:44] > in_mem[7][47:44]) begin
			in_mem[7][47:44] <= r2_data[7][47:44];
		end
		else begin
			in_mem[7][47:44] <= in_mem[7][47:44];
		end

		if (r2_data[7][51:48] > in_mem[7][51:48]) begin
			in_mem[7][51:48] <= r2_data[7][51:48];
		end
		else begin
			in_mem[7][51:48] <= in_mem[7][51:48];
		end

		if (r2_data[7][55:52] > in_mem[7][55:52]) begin
			in_mem[7][55:52] <= r2_data[7][55:52];
		end
		else begin
			in_mem[7][55:52] <= in_mem[7][55:52];
		end

		if (r2_data[7][59:56] > in_mem[7][59:56]) begin
			in_mem[7][59:56] <= r2_data[7][59:56];
		end
		else begin
			in_mem[7][59:56] <= in_mem[7][59:56];
		end

		if (r2_data[7][63:60] > in_mem[7][63:60]) begin
			in_mem[7][63:60] <= r2_data[7][63:60];
		end
		else begin
			in_mem[7][63:60] <= in_mem[7][63:60];
		end
	end
	else begin

		if (r2_data[7][3:0] > out_mem[7][3:0]) begin
			in_mem[7][3:0] <= r2_data[7][3:0];
		end
		else begin
			in_mem[7][3:0] <= out_mem[7][3:0];
		end

		if (r2_data[7][7:4] > out_mem[7][7:4]) begin
			in_mem[7][7:4] <= r2_data[7][7:4];
		end
		else begin
			in_mem[7][7:4] <= out_mem[7][7:4];
		end

		if (r2_data[7][11:8] > out_mem[7][11:8]) begin
			in_mem[7][11:8] <= r2_data[7][11:8];
		end
		else begin
			in_mem[7][11:8] <= out_mem[7][11:8];
		end

		if (r2_data[7][15:12] > out_mem[7][15:12]) begin
			in_mem[7][15:12] <= r2_data[7][15:12];
		end
		else begin
			in_mem[7][15:12] <= out_mem[7][15:12];
		end

		if (r2_data[7][19:16] > out_mem[7][19:16]) begin
			in_mem[7][19:16] <= r2_data[7][19:16];
		end
		else begin
			in_mem[7][19:16] <= out_mem[7][19:16];
		end

		if (r2_data[7][23:20] > out_mem[7][23:20]) begin
			in_mem[7][23:20] <= r2_data[7][23:20];
		end
		else begin
			in_mem[7][23:20] <= out_mem[7][23:20];
		end

		if (r2_data[7][27:24] > out_mem[7][27:24]) begin
			in_mem[7][27:24] <= r2_data[7][27:24];
		end
		else begin
			in_mem[7][27:24] <= out_mem[7][27:24];
		end

		if (r2_data[7][31:28] > out_mem[7][31:28]) begin
			in_mem[7][31:28] <= r2_data[7][31:28];
		end
		else begin
			in_mem[7][31:28] <= out_mem[7][31:28];
		end

		if (r2_data[7][35:32] > out_mem[7][35:32]) begin
			in_mem[7][35:32] <= r2_data[7][35:32];
		end
		else begin
			in_mem[7][35:32] <= out_mem[7][35:32];
		end

		if (r2_data[7][39:36] > out_mem[7][39:36]) begin
			in_mem[7][39:36] <= r2_data[7][39:36];
		end
		else begin
			in_mem[7][39:36] <= out_mem[7][39:36];
		end

		if (r2_data[7][43:40] > out_mem[7][43:40]) begin
			in_mem[7][43:40] <= r2_data[7][43:40];
		end
		else begin
			in_mem[7][43:40] <= out_mem[7][43:40];
		end

		if (r2_data[7][47:44] > out_mem[7][47:44]) begin
			in_mem[7][47:44] <= r2_data[7][47:44];
		end
		else begin
			in_mem[7][47:44] <= out_mem[7][47:44];
		end

		if (r2_data[7][51:48] > out_mem[7][51:48]) begin
			in_mem[7][51:48] <= r2_data[7][51:48];
		end
		else begin
			in_mem[7][51:48] <= out_mem[7][51:48];
		end

		if (r2_data[7][55:52] > out_mem[7][55:52]) begin
			in_mem[7][55:52] <= r2_data[7][55:52];
		end
		else begin
			in_mem[7][55:52] <= out_mem[7][55:52];
		end

		if (r2_data[7][59:56] > out_mem[7][59:56]) begin
			in_mem[7][59:56] <= r2_data[7][59:56];
		end
		else begin
			in_mem[7][59:56] <= out_mem[7][59:56];
		end

		if (r2_data[7][63:60] > out_mem[7][63:60]) begin
			in_mem[7][63:60] <= r2_data[7][63:60];
		end
		else begin
			in_mem[7][63:60] <= out_mem[7][63:60];
		end
	end
end

always_ff @(posedge clk) begin
	out_mem_valid <= {out_mem_valid, reading_memory};
	out_valid_in <= out_mem_valid[3];
	out_data_in <= max_tree_2[0];

	if (out_mem[0][3:0] > out_mem[1][3:0]) begin
		max_tree_0[0][3:0] <= out_mem[0][3:0];
	end
	else begin
		max_tree_0[0][3:0] <= out_mem[1][3:0];
	end

	if (out_mem[0][7:4] > out_mem[1][7:4]) begin
		max_tree_0[0][7:4] <= out_mem[0][7:4];
	end
	else begin
		max_tree_0[0][7:4] <= out_mem[1][7:4];
	end

	if (out_mem[0][11:8] > out_mem[1][11:8]) begin
		max_tree_0[0][11:8] <= out_mem[0][11:8];
	end
	else begin
		max_tree_0[0][11:8] <= out_mem[1][11:8];
	end

	if (out_mem[0][15:12] > out_mem[1][15:12]) begin
		max_tree_0[0][15:12] <= out_mem[0][15:12];
	end
	else begin
		max_tree_0[0][15:12] <= out_mem[1][15:12];
	end

	if (out_mem[0][19:16] > out_mem[1][19:16]) begin
		max_tree_0[0][19:16] <= out_mem[0][19:16];
	end
	else begin
		max_tree_0[0][19:16] <= out_mem[1][19:16];
	end

	if (out_mem[0][23:20] > out_mem[1][23:20]) begin
		max_tree_0[0][23:20] <= out_mem[0][23:20];
	end
	else begin
		max_tree_0[0][23:20] <= out_mem[1][23:20];
	end

	if (out_mem[0][27:24] > out_mem[1][27:24]) begin
		max_tree_0[0][27:24] <= out_mem[0][27:24];
	end
	else begin
		max_tree_0[0][27:24] <= out_mem[1][27:24];
	end

	if (out_mem[0][31:28] > out_mem[1][31:28]) begin
		max_tree_0[0][31:28] <= out_mem[0][31:28];
	end
	else begin
		max_tree_0[0][31:28] <= out_mem[1][31:28];
	end

	if (out_mem[0][35:32] > out_mem[1][35:32]) begin
		max_tree_0[0][35:32] <= out_mem[0][35:32];
	end
	else begin
		max_tree_0[0][35:32] <= out_mem[1][35:32];
	end

	if (out_mem[0][39:36] > out_mem[1][39:36]) begin
		max_tree_0[0][39:36] <= out_mem[0][39:36];
	end
	else begin
		max_tree_0[0][39:36] <= out_mem[1][39:36];
	end

	if (out_mem[0][43:40] > out_mem[1][43:40]) begin
		max_tree_0[0][43:40] <= out_mem[0][43:40];
	end
	else begin
		max_tree_0[0][43:40] <= out_mem[1][43:40];
	end

	if (out_mem[0][47:44] > out_mem[1][47:44]) begin
		max_tree_0[0][47:44] <= out_mem[0][47:44];
	end
	else begin
		max_tree_0[0][47:44] <= out_mem[1][47:44];
	end

	if (out_mem[0][51:48] > out_mem[1][51:48]) begin
		max_tree_0[0][51:48] <= out_mem[0][51:48];
	end
	else begin
		max_tree_0[0][51:48] <= out_mem[1][51:48];
	end

	if (out_mem[0][55:52] > out_mem[1][55:52]) begin
		max_tree_0[0][55:52] <= out_mem[0][55:52];
	end
	else begin
		max_tree_0[0][55:52] <= out_mem[1][55:52];
	end

	if (out_mem[0][59:56] > out_mem[1][59:56]) begin
		max_tree_0[0][59:56] <= out_mem[0][59:56];
	end
	else begin
		max_tree_0[0][59:56] <= out_mem[1][59:56];
	end

	if (out_mem[0][63:60] > out_mem[1][63:60]) begin
		max_tree_0[0][63:60] <= out_mem[0][63:60];
	end
	else begin
		max_tree_0[0][63:60] <= out_mem[1][63:60];
	end

	if (out_mem[2][3:0] > out_mem[3][3:0]) begin
		max_tree_0[1][3:0] <= out_mem[2][3:0];
	end
	else begin
		max_tree_0[1][3:0] <= out_mem[3][3:0];
	end

	if (out_mem[2][7:4] > out_mem[3][7:4]) begin
		max_tree_0[1][7:4] <= out_mem[2][7:4];
	end
	else begin
		max_tree_0[1][7:4] <= out_mem[3][7:4];
	end

	if (out_mem[2][11:8] > out_mem[3][11:8]) begin
		max_tree_0[1][11:8] <= out_mem[2][11:8];
	end
	else begin
		max_tree_0[1][11:8] <= out_mem[3][11:8];
	end

	if (out_mem[2][15:12] > out_mem[3][15:12]) begin
		max_tree_0[1][15:12] <= out_mem[2][15:12];
	end
	else begin
		max_tree_0[1][15:12] <= out_mem[3][15:12];
	end

	if (out_mem[2][19:16] > out_mem[3][19:16]) begin
		max_tree_0[1][19:16] <= out_mem[2][19:16];
	end
	else begin
		max_tree_0[1][19:16] <= out_mem[3][19:16];
	end

	if (out_mem[2][23:20] > out_mem[3][23:20]) begin
		max_tree_0[1][23:20] <= out_mem[2][23:20];
	end
	else begin
		max_tree_0[1][23:20] <= out_mem[3][23:20];
	end

	if (out_mem[2][27:24] > out_mem[3][27:24]) begin
		max_tree_0[1][27:24] <= out_mem[2][27:24];
	end
	else begin
		max_tree_0[1][27:24] <= out_mem[3][27:24];
	end

	if (out_mem[2][31:28] > out_mem[3][31:28]) begin
		max_tree_0[1][31:28] <= out_mem[2][31:28];
	end
	else begin
		max_tree_0[1][31:28] <= out_mem[3][31:28];
	end

	if (out_mem[2][35:32] > out_mem[3][35:32]) begin
		max_tree_0[1][35:32] <= out_mem[2][35:32];
	end
	else begin
		max_tree_0[1][35:32] <= out_mem[3][35:32];
	end

	if (out_mem[2][39:36] > out_mem[3][39:36]) begin
		max_tree_0[1][39:36] <= out_mem[2][39:36];
	end
	else begin
		max_tree_0[1][39:36] <= out_mem[3][39:36];
	end

	if (out_mem[2][43:40] > out_mem[3][43:40]) begin
		max_tree_0[1][43:40] <= out_mem[2][43:40];
	end
	else begin
		max_tree_0[1][43:40] <= out_mem[3][43:40];
	end

	if (out_mem[2][47:44] > out_mem[3][47:44]) begin
		max_tree_0[1][47:44] <= out_mem[2][47:44];
	end
	else begin
		max_tree_0[1][47:44] <= out_mem[3][47:44];
	end

	if (out_mem[2][51:48] > out_mem[3][51:48]) begin
		max_tree_0[1][51:48] <= out_mem[2][51:48];
	end
	else begin
		max_tree_0[1][51:48] <= out_mem[3][51:48];
	end

	if (out_mem[2][55:52] > out_mem[3][55:52]) begin
		max_tree_0[1][55:52] <= out_mem[2][55:52];
	end
	else begin
		max_tree_0[1][55:52] <= out_mem[3][55:52];
	end

	if (out_mem[2][59:56] > out_mem[3][59:56]) begin
		max_tree_0[1][59:56] <= out_mem[2][59:56];
	end
	else begin
		max_tree_0[1][59:56] <= out_mem[3][59:56];
	end

	if (out_mem[2][63:60] > out_mem[3][63:60]) begin
		max_tree_0[1][63:60] <= out_mem[2][63:60];
	end
	else begin
		max_tree_0[1][63:60] <= out_mem[3][63:60];
	end

	if (out_mem[4][3:0] > out_mem[5][3:0]) begin
		max_tree_0[2][3:0] <= out_mem[4][3:0];
	end
	else begin
		max_tree_0[2][3:0] <= out_mem[5][3:0];
	end

	if (out_mem[4][7:4] > out_mem[5][7:4]) begin
		max_tree_0[2][7:4] <= out_mem[4][7:4];
	end
	else begin
		max_tree_0[2][7:4] <= out_mem[5][7:4];
	end

	if (out_mem[4][11:8] > out_mem[5][11:8]) begin
		max_tree_0[2][11:8] <= out_mem[4][11:8];
	end
	else begin
		max_tree_0[2][11:8] <= out_mem[5][11:8];
	end

	if (out_mem[4][15:12] > out_mem[5][15:12]) begin
		max_tree_0[2][15:12] <= out_mem[4][15:12];
	end
	else begin
		max_tree_0[2][15:12] <= out_mem[5][15:12];
	end

	if (out_mem[4][19:16] > out_mem[5][19:16]) begin
		max_tree_0[2][19:16] <= out_mem[4][19:16];
	end
	else begin
		max_tree_0[2][19:16] <= out_mem[5][19:16];
	end

	if (out_mem[4][23:20] > out_mem[5][23:20]) begin
		max_tree_0[2][23:20] <= out_mem[4][23:20];
	end
	else begin
		max_tree_0[2][23:20] <= out_mem[5][23:20];
	end

	if (out_mem[4][27:24] > out_mem[5][27:24]) begin
		max_tree_0[2][27:24] <= out_mem[4][27:24];
	end
	else begin
		max_tree_0[2][27:24] <= out_mem[5][27:24];
	end

	if (out_mem[4][31:28] > out_mem[5][31:28]) begin
		max_tree_0[2][31:28] <= out_mem[4][31:28];
	end
	else begin
		max_tree_0[2][31:28] <= out_mem[5][31:28];
	end

	if (out_mem[4][35:32] > out_mem[5][35:32]) begin
		max_tree_0[2][35:32] <= out_mem[4][35:32];
	end
	else begin
		max_tree_0[2][35:32] <= out_mem[5][35:32];
	end

	if (out_mem[4][39:36] > out_mem[5][39:36]) begin
		max_tree_0[2][39:36] <= out_mem[4][39:36];
	end
	else begin
		max_tree_0[2][39:36] <= out_mem[5][39:36];
	end

	if (out_mem[4][43:40] > out_mem[5][43:40]) begin
		max_tree_0[2][43:40] <= out_mem[4][43:40];
	end
	else begin
		max_tree_0[2][43:40] <= out_mem[5][43:40];
	end

	if (out_mem[4][47:44] > out_mem[5][47:44]) begin
		max_tree_0[2][47:44] <= out_mem[4][47:44];
	end
	else begin
		max_tree_0[2][47:44] <= out_mem[5][47:44];
	end

	if (out_mem[4][51:48] > out_mem[5][51:48]) begin
		max_tree_0[2][51:48] <= out_mem[4][51:48];
	end
	else begin
		max_tree_0[2][51:48] <= out_mem[5][51:48];
	end

	if (out_mem[4][55:52] > out_mem[5][55:52]) begin
		max_tree_0[2][55:52] <= out_mem[4][55:52];
	end
	else begin
		max_tree_0[2][55:52] <= out_mem[5][55:52];
	end

	if (out_mem[4][59:56] > out_mem[5][59:56]) begin
		max_tree_0[2][59:56] <= out_mem[4][59:56];
	end
	else begin
		max_tree_0[2][59:56] <= out_mem[5][59:56];
	end

	if (out_mem[4][63:60] > out_mem[5][63:60]) begin
		max_tree_0[2][63:60] <= out_mem[4][63:60];
	end
	else begin
		max_tree_0[2][63:60] <= out_mem[5][63:60];
	end

	if (out_mem[6][3:0] > out_mem[7][3:0]) begin
		max_tree_0[3][3:0] <= out_mem[6][3:0];
	end
	else begin
		max_tree_0[3][3:0] <= out_mem[7][3:0];
	end

	if (out_mem[6][7:4] > out_mem[7][7:4]) begin
		max_tree_0[3][7:4] <= out_mem[6][7:4];
	end
	else begin
		max_tree_0[3][7:4] <= out_mem[7][7:4];
	end

	if (out_mem[6][11:8] > out_mem[7][11:8]) begin
		max_tree_0[3][11:8] <= out_mem[6][11:8];
	end
	else begin
		max_tree_0[3][11:8] <= out_mem[7][11:8];
	end

	if (out_mem[6][15:12] > out_mem[7][15:12]) begin
		max_tree_0[3][15:12] <= out_mem[6][15:12];
	end
	else begin
		max_tree_0[3][15:12] <= out_mem[7][15:12];
	end

	if (out_mem[6][19:16] > out_mem[7][19:16]) begin
		max_tree_0[3][19:16] <= out_mem[6][19:16];
	end
	else begin
		max_tree_0[3][19:16] <= out_mem[7][19:16];
	end

	if (out_mem[6][23:20] > out_mem[7][23:20]) begin
		max_tree_0[3][23:20] <= out_mem[6][23:20];
	end
	else begin
		max_tree_0[3][23:20] <= out_mem[7][23:20];
	end

	if (out_mem[6][27:24] > out_mem[7][27:24]) begin
		max_tree_0[3][27:24] <= out_mem[6][27:24];
	end
	else begin
		max_tree_0[3][27:24] <= out_mem[7][27:24];
	end

	if (out_mem[6][31:28] > out_mem[7][31:28]) begin
		max_tree_0[3][31:28] <= out_mem[6][31:28];
	end
	else begin
		max_tree_0[3][31:28] <= out_mem[7][31:28];
	end

	if (out_mem[6][35:32] > out_mem[7][35:32]) begin
		max_tree_0[3][35:32] <= out_mem[6][35:32];
	end
	else begin
		max_tree_0[3][35:32] <= out_mem[7][35:32];
	end

	if (out_mem[6][39:36] > out_mem[7][39:36]) begin
		max_tree_0[3][39:36] <= out_mem[6][39:36];
	end
	else begin
		max_tree_0[3][39:36] <= out_mem[7][39:36];
	end

	if (out_mem[6][43:40] > out_mem[7][43:40]) begin
		max_tree_0[3][43:40] <= out_mem[6][43:40];
	end
	else begin
		max_tree_0[3][43:40] <= out_mem[7][43:40];
	end

	if (out_mem[6][47:44] > out_mem[7][47:44]) begin
		max_tree_0[3][47:44] <= out_mem[6][47:44];
	end
	else begin
		max_tree_0[3][47:44] <= out_mem[7][47:44];
	end

	if (out_mem[6][51:48] > out_mem[7][51:48]) begin
		max_tree_0[3][51:48] <= out_mem[6][51:48];
	end
	else begin
		max_tree_0[3][51:48] <= out_mem[7][51:48];
	end

	if (out_mem[6][55:52] > out_mem[7][55:52]) begin
		max_tree_0[3][55:52] <= out_mem[6][55:52];
	end
	else begin
		max_tree_0[3][55:52] <= out_mem[7][55:52];
	end

	if (out_mem[6][59:56] > out_mem[7][59:56]) begin
		max_tree_0[3][59:56] <= out_mem[6][59:56];
	end
	else begin
		max_tree_0[3][59:56] <= out_mem[7][59:56];
	end

	if (out_mem[6][63:60] > out_mem[7][63:60]) begin
		max_tree_0[3][63:60] <= out_mem[6][63:60];
	end
	else begin
		max_tree_0[3][63:60] <= out_mem[7][63:60];
	end

	if (max_tree_0[0][3:0] > max_tree_0[1][3:0]) begin
		max_tree_1[0][3:0] <= max_tree_0[0][3:0];
	end
	else begin
		max_tree_1[0][3:0] <= max_tree_0[1][3:0];
	end

	if (max_tree_0[0][7:4] > max_tree_0[1][7:4]) begin
		max_tree_1[0][7:4] <= max_tree_0[0][7:4];
	end
	else begin
		max_tree_1[0][7:4] <= max_tree_0[1][7:4];
	end

	if (max_tree_0[0][11:8] > max_tree_0[1][11:8]) begin
		max_tree_1[0][11:8] <= max_tree_0[0][11:8];
	end
	else begin
		max_tree_1[0][11:8] <= max_tree_0[1][11:8];
	end

	if (max_tree_0[0][15:12] > max_tree_0[1][15:12]) begin
		max_tree_1[0][15:12] <= max_tree_0[0][15:12];
	end
	else begin
		max_tree_1[0][15:12] <= max_tree_0[1][15:12];
	end

	if (max_tree_0[0][19:16] > max_tree_0[1][19:16]) begin
		max_tree_1[0][19:16] <= max_tree_0[0][19:16];
	end
	else begin
		max_tree_1[0][19:16] <= max_tree_0[1][19:16];
	end

	if (max_tree_0[0][23:20] > max_tree_0[1][23:20]) begin
		max_tree_1[0][23:20] <= max_tree_0[0][23:20];
	end
	else begin
		max_tree_1[0][23:20] <= max_tree_0[1][23:20];
	end

	if (max_tree_0[0][27:24] > max_tree_0[1][27:24]) begin
		max_tree_1[0][27:24] <= max_tree_0[0][27:24];
	end
	else begin
		max_tree_1[0][27:24] <= max_tree_0[1][27:24];
	end

	if (max_tree_0[0][31:28] > max_tree_0[1][31:28]) begin
		max_tree_1[0][31:28] <= max_tree_0[0][31:28];
	end
	else begin
		max_tree_1[0][31:28] <= max_tree_0[1][31:28];
	end

	if (max_tree_0[0][35:32] > max_tree_0[1][35:32]) begin
		max_tree_1[0][35:32] <= max_tree_0[0][35:32];
	end
	else begin
		max_tree_1[0][35:32] <= max_tree_0[1][35:32];
	end

	if (max_tree_0[0][39:36] > max_tree_0[1][39:36]) begin
		max_tree_1[0][39:36] <= max_tree_0[0][39:36];
	end
	else begin
		max_tree_1[0][39:36] <= max_tree_0[1][39:36];
	end

	if (max_tree_0[0][43:40] > max_tree_0[1][43:40]) begin
		max_tree_1[0][43:40] <= max_tree_0[0][43:40];
	end
	else begin
		max_tree_1[0][43:40] <= max_tree_0[1][43:40];
	end

	if (max_tree_0[0][47:44] > max_tree_0[1][47:44]) begin
		max_tree_1[0][47:44] <= max_tree_0[0][47:44];
	end
	else begin
		max_tree_1[0][47:44] <= max_tree_0[1][47:44];
	end

	if (max_tree_0[0][51:48] > max_tree_0[1][51:48]) begin
		max_tree_1[0][51:48] <= max_tree_0[0][51:48];
	end
	else begin
		max_tree_1[0][51:48] <= max_tree_0[1][51:48];
	end

	if (max_tree_0[0][55:52] > max_tree_0[1][55:52]) begin
		max_tree_1[0][55:52] <= max_tree_0[0][55:52];
	end
	else begin
		max_tree_1[0][55:52] <= max_tree_0[1][55:52];
	end

	if (max_tree_0[0][59:56] > max_tree_0[1][59:56]) begin
		max_tree_1[0][59:56] <= max_tree_0[0][59:56];
	end
	else begin
		max_tree_1[0][59:56] <= max_tree_0[1][59:56];
	end

	if (max_tree_0[0][63:60] > max_tree_0[1][63:60]) begin
		max_tree_1[0][63:60] <= max_tree_0[0][63:60];
	end
	else begin
		max_tree_1[0][63:60] <= max_tree_0[1][63:60];
	end

	if (max_tree_0[2][3:0] > max_tree_0[3][3:0]) begin
		max_tree_1[1][3:0] <= max_tree_0[2][3:0];
	end
	else begin
		max_tree_1[1][3:0] <= max_tree_0[3][3:0];
	end

	if (max_tree_0[2][7:4] > max_tree_0[3][7:4]) begin
		max_tree_1[1][7:4] <= max_tree_0[2][7:4];
	end
	else begin
		max_tree_1[1][7:4] <= max_tree_0[3][7:4];
	end

	if (max_tree_0[2][11:8] > max_tree_0[3][11:8]) begin
		max_tree_1[1][11:8] <= max_tree_0[2][11:8];
	end
	else begin
		max_tree_1[1][11:8] <= max_tree_0[3][11:8];
	end

	if (max_tree_0[2][15:12] > max_tree_0[3][15:12]) begin
		max_tree_1[1][15:12] <= max_tree_0[2][15:12];
	end
	else begin
		max_tree_1[1][15:12] <= max_tree_0[3][15:12];
	end

	if (max_tree_0[2][19:16] > max_tree_0[3][19:16]) begin
		max_tree_1[1][19:16] <= max_tree_0[2][19:16];
	end
	else begin
		max_tree_1[1][19:16] <= max_tree_0[3][19:16];
	end

	if (max_tree_0[2][23:20] > max_tree_0[3][23:20]) begin
		max_tree_1[1][23:20] <= max_tree_0[2][23:20];
	end
	else begin
		max_tree_1[1][23:20] <= max_tree_0[3][23:20];
	end

	if (max_tree_0[2][27:24] > max_tree_0[3][27:24]) begin
		max_tree_1[1][27:24] <= max_tree_0[2][27:24];
	end
	else begin
		max_tree_1[1][27:24] <= max_tree_0[3][27:24];
	end

	if (max_tree_0[2][31:28] > max_tree_0[3][31:28]) begin
		max_tree_1[1][31:28] <= max_tree_0[2][31:28];
	end
	else begin
		max_tree_1[1][31:28] <= max_tree_0[3][31:28];
	end

	if (max_tree_0[2][35:32] > max_tree_0[3][35:32]) begin
		max_tree_1[1][35:32] <= max_tree_0[2][35:32];
	end
	else begin
		max_tree_1[1][35:32] <= max_tree_0[3][35:32];
	end

	if (max_tree_0[2][39:36] > max_tree_0[3][39:36]) begin
		max_tree_1[1][39:36] <= max_tree_0[2][39:36];
	end
	else begin
		max_tree_1[1][39:36] <= max_tree_0[3][39:36];
	end

	if (max_tree_0[2][43:40] > max_tree_0[3][43:40]) begin
		max_tree_1[1][43:40] <= max_tree_0[2][43:40];
	end
	else begin
		max_tree_1[1][43:40] <= max_tree_0[3][43:40];
	end

	if (max_tree_0[2][47:44] > max_tree_0[3][47:44]) begin
		max_tree_1[1][47:44] <= max_tree_0[2][47:44];
	end
	else begin
		max_tree_1[1][47:44] <= max_tree_0[3][47:44];
	end

	if (max_tree_0[2][51:48] > max_tree_0[3][51:48]) begin
		max_tree_1[1][51:48] <= max_tree_0[2][51:48];
	end
	else begin
		max_tree_1[1][51:48] <= max_tree_0[3][51:48];
	end

	if (max_tree_0[2][55:52] > max_tree_0[3][55:52]) begin
		max_tree_1[1][55:52] <= max_tree_0[2][55:52];
	end
	else begin
		max_tree_1[1][55:52] <= max_tree_0[3][55:52];
	end

	if (max_tree_0[2][59:56] > max_tree_0[3][59:56]) begin
		max_tree_1[1][59:56] <= max_tree_0[2][59:56];
	end
	else begin
		max_tree_1[1][59:56] <= max_tree_0[3][59:56];
	end

	if (max_tree_0[2][63:60] > max_tree_0[3][63:60]) begin
		max_tree_1[1][63:60] <= max_tree_0[2][63:60];
	end
	else begin
		max_tree_1[1][63:60] <= max_tree_0[3][63:60];
	end

	if (max_tree_1[0][3:0] > max_tree_1[1][3:0]) begin
		max_tree_2[0][3:0] <= max_tree_1[0][3:0];
	end
	else begin
		max_tree_2[0][3:0] <= max_tree_1[1][3:0];
	end

	if (max_tree_1[0][7:4] > max_tree_1[1][7:4]) begin
		max_tree_2[0][7:4] <= max_tree_1[0][7:4];
	end
	else begin
		max_tree_2[0][7:4] <= max_tree_1[1][7:4];
	end

	if (max_tree_1[0][11:8] > max_tree_1[1][11:8]) begin
		max_tree_2[0][11:8] <= max_tree_1[0][11:8];
	end
	else begin
		max_tree_2[0][11:8] <= max_tree_1[1][11:8];
	end

	if (max_tree_1[0][15:12] > max_tree_1[1][15:12]) begin
		max_tree_2[0][15:12] <= max_tree_1[0][15:12];
	end
	else begin
		max_tree_2[0][15:12] <= max_tree_1[1][15:12];
	end

	if (max_tree_1[0][19:16] > max_tree_1[1][19:16]) begin
		max_tree_2[0][19:16] <= max_tree_1[0][19:16];
	end
	else begin
		max_tree_2[0][19:16] <= max_tree_1[1][19:16];
	end

	if (max_tree_1[0][23:20] > max_tree_1[1][23:20]) begin
		max_tree_2[0][23:20] <= max_tree_1[0][23:20];
	end
	else begin
		max_tree_2[0][23:20] <= max_tree_1[1][23:20];
	end

	if (max_tree_1[0][27:24] > max_tree_1[1][27:24]) begin
		max_tree_2[0][27:24] <= max_tree_1[0][27:24];
	end
	else begin
		max_tree_2[0][27:24] <= max_tree_1[1][27:24];
	end

	if (max_tree_1[0][31:28] > max_tree_1[1][31:28]) begin
		max_tree_2[0][31:28] <= max_tree_1[0][31:28];
	end
	else begin
		max_tree_2[0][31:28] <= max_tree_1[1][31:28];
	end

	if (max_tree_1[0][35:32] > max_tree_1[1][35:32]) begin
		max_tree_2[0][35:32] <= max_tree_1[0][35:32];
	end
	else begin
		max_tree_2[0][35:32] <= max_tree_1[1][35:32];
	end

	if (max_tree_1[0][39:36] > max_tree_1[1][39:36]) begin
		max_tree_2[0][39:36] <= max_tree_1[0][39:36];
	end
	else begin
		max_tree_2[0][39:36] <= max_tree_1[1][39:36];
	end

	if (max_tree_1[0][43:40] > max_tree_1[1][43:40]) begin
		max_tree_2[0][43:40] <= max_tree_1[0][43:40];
	end
	else begin
		max_tree_2[0][43:40] <= max_tree_1[1][43:40];
	end

	if (max_tree_1[0][47:44] > max_tree_1[1][47:44]) begin
		max_tree_2[0][47:44] <= max_tree_1[0][47:44];
	end
	else begin
		max_tree_2[0][47:44] <= max_tree_1[1][47:44];
	end

	if (max_tree_1[0][51:48] > max_tree_1[1][51:48]) begin
		max_tree_2[0][51:48] <= max_tree_1[0][51:48];
	end
	else begin
		max_tree_2[0][51:48] <= max_tree_1[1][51:48];
	end

	if (max_tree_1[0][55:52] > max_tree_1[1][55:52]) begin
		max_tree_2[0][55:52] <= max_tree_1[0][55:52];
	end
	else begin
		max_tree_2[0][55:52] <= max_tree_1[1][55:52];
	end

	if (max_tree_1[0][59:56] > max_tree_1[1][59:56]) begin
		max_tree_2[0][59:56] <= max_tree_1[0][59:56];
	end
	else begin
		max_tree_2[0][59:56] <= max_tree_1[1][59:56];
	end

	if (max_tree_1[0][63:60] > max_tree_1[1][63:60]) begin
		max_tree_2[0][63:60] <= max_tree_1[0][63:60];
	end
	else begin
		max_tree_2[0][63:60] <= max_tree_1[1][63:60];
	end
end

always_ff @(posedge clk) begin
	out_data <= {out_data_in, out_data[511:64]};

	if (out_valid_in) begin

		if (out_valid_cnt == 4'd7) begin
			out_valid_cnt <= 4'd0;
			out_valid <= out_ready;
		end
		else begin
			out_valid_cnt <= out_valid_cnt + 4'd1;
			out_valid <= 1'd0;
		end
	end
	else begin
		out_valid_cnt <= out_valid_cnt;
		out_valid <= 1'd0;
	end
end

endmodule

